library ieee;
use ieee.std_logic_1164.all;
-- Uncomment the following line if VHDL primitives are in use.
-- use prims.all;
entity rwcomp0 is
  Port ( clk : in std_logic ;
         input : in std_logic_vector (0 to 639);
         output : out std_logic_vector (0 to 511));
end rwcomp0;

architecture behavioral of rwcomp0 is
  type control_state is (STATE0,STATE1163,STATE3537);
  function rewire_key2_3233 return std_logic_vector;
  function rewire_key1_2939 return std_logic_vector;
  function rewire_buildSalsa256_1182(r1183 : std_logic_vector ; r1184 : std_logic_vector ; r1185 : std_logic_vector ; r1186 : std_logic_vector) return std_logic_vector;
  function rewire_salsaHash_1658(r1659 : std_logic_vector) return std_logic_vector;
  function rewire_impwords_2602(r2603 : std_logic_vector) return std_logic_vector;
  function rewire_littleendian_2736(r2737 : std_logic_vector) return std_logic_vector;
  function rewire_w8to16le_2831(r2832 : std_logic_vector ; r2833 : std_logic_vector) return std_logic_vector;
  function rewire_w16tow32le_2750(r2751 : std_logic_vector ; r2752 : std_logic_vector) return std_logic_vector;
  function rewire_salsaHashp_1978(r1979 : std_logic_vector) return std_logic_vector;
  function rewire_doubleRound_2016(r2017 : std_logic_vector) return std_logic_vector;
  function rewire_columnRound_2436(r2437 : std_logic_vector) return std_logic_vector;
  function rewire_rowRound_2019(r2020 : std_logic_vector) return std_logic_vector;
  function rewire_quarterRound_2057(r2058 : std_logic_vector) return std_logic_vector;
  function rewire_rot18_2296(r2297 : std_logic_vector) return std_logic_vector;
  function rewire_rot13_2221(r2222 : std_logic_vector) return std_logic_vector;
  function rewire_rot9_2146(r2147 : std_logic_vector) return std_logic_vector;
  function rewire_rot7_2071(r2072 : std_logic_vector) return std_logic_vector;
  function rewire_expwords_1661(r1662 : std_logic_vector) return std_logic_vector;
  function rewire_littleendianp_1699(r1700 : std_logic_vector) return std_logic_vector;
  function rewire_sigma3_1533 return std_logic_vector;
  function rewire_sigma2_1456 return std_logic_vector;
  function rewire_sigma1_1379 return std_logic_vector;
  function rewire_sigma0_1302 return std_logic_vector;
  function rewire_zerothoutput_3 return std_logic_vector;

  function rewire_key2_3233 return std_logic_vector
  is
    variable r3524 : std_logic_vector(0 to 127) := (others => '0');
    variable r3523 : std_logic_vector(0 to 7) := (others => '0');
    variable r3521 : std_logic_vector(0 to 0) := (others => '0');
    variable r3519 : std_logic_vector(0 to 0) := (others => '0');
    variable r3517 : std_logic_vector(0 to 0) := (others => '0');
    variable r3515 : std_logic_vector(0 to 0) := (others => '0');
    variable r3513 : std_logic_vector(0 to 0) := (others => '0');
    variable r3511 : std_logic_vector(0 to 0) := (others => '0');
    variable r3509 : std_logic_vector(0 to 0) := (others => '0');
    variable r3507 : std_logic_vector(0 to 0) := (others => '0');
    variable r3505 : std_logic_vector(0 to 7) := (others => '0');
    variable r3503 : std_logic_vector(0 to 0) := (others => '0');
    variable r3501 : std_logic_vector(0 to 0) := (others => '0');
    variable r3499 : std_logic_vector(0 to 0) := (others => '0');
    variable r3497 : std_logic_vector(0 to 0) := (others => '0');
    variable r3495 : std_logic_vector(0 to 0) := (others => '0');
    variable r3493 : std_logic_vector(0 to 0) := (others => '0');
    variable r3491 : std_logic_vector(0 to 0) := (others => '0');
    variable r3489 : std_logic_vector(0 to 0) := (others => '0');
    variable r3487 : std_logic_vector(0 to 7) := (others => '0');
    variable r3485 : std_logic_vector(0 to 0) := (others => '0');
    variable r3483 : std_logic_vector(0 to 0) := (others => '0');
    variable r3481 : std_logic_vector(0 to 0) := (others => '0');
    variable r3479 : std_logic_vector(0 to 0) := (others => '0');
    variable r3477 : std_logic_vector(0 to 0) := (others => '0');
    variable r3475 : std_logic_vector(0 to 0) := (others => '0');
    variable r3473 : std_logic_vector(0 to 0) := (others => '0');
    variable r3471 : std_logic_vector(0 to 0) := (others => '0');
    variable r3469 : std_logic_vector(0 to 7) := (others => '0');
    variable r3467 : std_logic_vector(0 to 0) := (others => '0');
    variable r3465 : std_logic_vector(0 to 0) := (others => '0');
    variable r3463 : std_logic_vector(0 to 0) := (others => '0');
    variable r3461 : std_logic_vector(0 to 0) := (others => '0');
    variable r3459 : std_logic_vector(0 to 0) := (others => '0');
    variable r3457 : std_logic_vector(0 to 0) := (others => '0');
    variable r3455 : std_logic_vector(0 to 0) := (others => '0');
    variable r3453 : std_logic_vector(0 to 0) := (others => '0');
    variable r3451 : std_logic_vector(0 to 7) := (others => '0');
    variable r3449 : std_logic_vector(0 to 0) := (others => '0');
    variable r3447 : std_logic_vector(0 to 0) := (others => '0');
    variable r3445 : std_logic_vector(0 to 0) := (others => '0');
    variable r3443 : std_logic_vector(0 to 0) := (others => '0');
    variable r3441 : std_logic_vector(0 to 0) := (others => '0');
    variable r3439 : std_logic_vector(0 to 0) := (others => '0');
    variable r3437 : std_logic_vector(0 to 0) := (others => '0');
    variable r3435 : std_logic_vector(0 to 0) := (others => '0');
    variable r3433 : std_logic_vector(0 to 7) := (others => '0');
    variable r3431 : std_logic_vector(0 to 0) := (others => '0');
    variable r3429 : std_logic_vector(0 to 0) := (others => '0');
    variable r3427 : std_logic_vector(0 to 0) := (others => '0');
    variable r3425 : std_logic_vector(0 to 0) := (others => '0');
    variable r3423 : std_logic_vector(0 to 0) := (others => '0');
    variable r3421 : std_logic_vector(0 to 0) := (others => '0');
    variable r3419 : std_logic_vector(0 to 0) := (others => '0');
    variable r3417 : std_logic_vector(0 to 0) := (others => '0');
    variable r3415 : std_logic_vector(0 to 7) := (others => '0');
    variable r3413 : std_logic_vector(0 to 0) := (others => '0');
    variable r3411 : std_logic_vector(0 to 0) := (others => '0');
    variable r3409 : std_logic_vector(0 to 0) := (others => '0');
    variable r3407 : std_logic_vector(0 to 0) := (others => '0');
    variable r3405 : std_logic_vector(0 to 0) := (others => '0');
    variable r3403 : std_logic_vector(0 to 0) := (others => '0');
    variable r3401 : std_logic_vector(0 to 0) := (others => '0');
    variable r3399 : std_logic_vector(0 to 0) := (others => '0');
    variable r3397 : std_logic_vector(0 to 7) := (others => '0');
    variable r3395 : std_logic_vector(0 to 0) := (others => '0');
    variable r3393 : std_logic_vector(0 to 0) := (others => '0');
    variable r3391 : std_logic_vector(0 to 0) := (others => '0');
    variable r3389 : std_logic_vector(0 to 0) := (others => '0');
    variable r3387 : std_logic_vector(0 to 0) := (others => '0');
    variable r3385 : std_logic_vector(0 to 0) := (others => '0');
    variable r3383 : std_logic_vector(0 to 0) := (others => '0');
    variable r3381 : std_logic_vector(0 to 0) := (others => '0');
    variable r3379 : std_logic_vector(0 to 7) := (others => '0');
    variable r3377 : std_logic_vector(0 to 0) := (others => '0');
    variable r3375 : std_logic_vector(0 to 0) := (others => '0');
    variable r3373 : std_logic_vector(0 to 0) := (others => '0');
    variable r3371 : std_logic_vector(0 to 0) := (others => '0');
    variable r3369 : std_logic_vector(0 to 0) := (others => '0');
    variable r3367 : std_logic_vector(0 to 0) := (others => '0');
    variable r3365 : std_logic_vector(0 to 0) := (others => '0');
    variable r3363 : std_logic_vector(0 to 0) := (others => '0');
    variable r3361 : std_logic_vector(0 to 7) := (others => '0');
    variable r3359 : std_logic_vector(0 to 0) := (others => '0');
    variable r3357 : std_logic_vector(0 to 0) := (others => '0');
    variable r3355 : std_logic_vector(0 to 0) := (others => '0');
    variable r3353 : std_logic_vector(0 to 0) := (others => '0');
    variable r3351 : std_logic_vector(0 to 0) := (others => '0');
    variable r3349 : std_logic_vector(0 to 0) := (others => '0');
    variable r3347 : std_logic_vector(0 to 0) := (others => '0');
    variable r3345 : std_logic_vector(0 to 0) := (others => '0');
    variable r3343 : std_logic_vector(0 to 7) := (others => '0');
    variable r3341 : std_logic_vector(0 to 0) := (others => '0');
    variable r3339 : std_logic_vector(0 to 0) := (others => '0');
    variable r3337 : std_logic_vector(0 to 0) := (others => '0');
    variable r3335 : std_logic_vector(0 to 0) := (others => '0');
    variable r3333 : std_logic_vector(0 to 0) := (others => '0');
    variable r3331 : std_logic_vector(0 to 0) := (others => '0');
    variable r3329 : std_logic_vector(0 to 0) := (others => '0');
    variable r3327 : std_logic_vector(0 to 0) := (others => '0');
    variable r3325 : std_logic_vector(0 to 7) := (others => '0');
    variable r3323 : std_logic_vector(0 to 0) := (others => '0');
    variable r3321 : std_logic_vector(0 to 0) := (others => '0');
    variable r3319 : std_logic_vector(0 to 0) := (others => '0');
    variable r3317 : std_logic_vector(0 to 0) := (others => '0');
    variable r3315 : std_logic_vector(0 to 0) := (others => '0');
    variable r3313 : std_logic_vector(0 to 0) := (others => '0');
    variable r3311 : std_logic_vector(0 to 0) := (others => '0');
    variable r3309 : std_logic_vector(0 to 0) := (others => '0');
    variable r3307 : std_logic_vector(0 to 7) := (others => '0');
    variable r3305 : std_logic_vector(0 to 0) := (others => '0');
    variable r3303 : std_logic_vector(0 to 0) := (others => '0');
    variable r3301 : std_logic_vector(0 to 0) := (others => '0');
    variable r3299 : std_logic_vector(0 to 0) := (others => '0');
    variable r3297 : std_logic_vector(0 to 0) := (others => '0');
    variable r3295 : std_logic_vector(0 to 0) := (others => '0');
    variable r3293 : std_logic_vector(0 to 0) := (others => '0');
    variable r3291 : std_logic_vector(0 to 0) := (others => '0');
    variable r3289 : std_logic_vector(0 to 7) := (others => '0');
    variable r3287 : std_logic_vector(0 to 0) := (others => '0');
    variable r3285 : std_logic_vector(0 to 0) := (others => '0');
    variable r3283 : std_logic_vector(0 to 0) := (others => '0');
    variable r3281 : std_logic_vector(0 to 0) := (others => '0');
    variable r3279 : std_logic_vector(0 to 0) := (others => '0');
    variable r3277 : std_logic_vector(0 to 0) := (others => '0');
    variable r3275 : std_logic_vector(0 to 0) := (others => '0');
    variable r3273 : std_logic_vector(0 to 0) := (others => '0');
    variable r3271 : std_logic_vector(0 to 7) := (others => '0');
    variable r3269 : std_logic_vector(0 to 0) := (others => '0');
    variable r3267 : std_logic_vector(0 to 0) := (others => '0');
    variable r3265 : std_logic_vector(0 to 0) := (others => '0');
    variable r3263 : std_logic_vector(0 to 0) := (others => '0');
    variable r3261 : std_logic_vector(0 to 0) := (others => '0');
    variable r3259 : std_logic_vector(0 to 0) := (others => '0');
    variable r3257 : std_logic_vector(0 to 0) := (others => '0');
    variable r3255 : std_logic_vector(0 to 0) := (others => '0');
    variable r3253 : std_logic_vector(0 to 7) := (others => '0');
    variable r3251 : std_logic_vector(0 to 0) := (others => '0');
    variable r3249 : std_logic_vector(0 to 0) := (others => '0');
    variable r3247 : std_logic_vector(0 to 0) := (others => '0');
    variable r3245 : std_logic_vector(0 to 0) := (others => '0');
    variable r3243 : std_logic_vector(0 to 0) := (others => '0');
    variable r3241 : std_logic_vector(0 to 0) := (others => '0');
    variable r3239 : std_logic_vector(0 to 0) := (others => '0');
    variable r3237 : std_logic_vector(0 to 0) := (others => '0');
  begin
    r3237 := "0";
    r3239 := "1";
    r3241 := "1";
    r3243 := "1";
    r3245 := "0";
    r3247 := "1";
    r3249 := "1";
    r3251 := "1";
    r3253 := (r3237 & r3239 & r3241 & r3243 & r3245 & r3247 & r3249 & r3251);
    r3255 := "1";
    r3257 := "0";
    r3259 := "1";
    r3261 := "1";
    r3263 := "0";
    r3265 := "1";
    r3267 := "1";
    r3269 := "1";
    r3271 := (r3255 & r3257 & r3259 & r3261 & r3263 & r3265 & r3267 & r3269);
    r3273 := "0";
    r3275 := "0";
    r3277 := "1";
    r3279 := "1";
    r3281 := "0";
    r3283 := "1";
    r3285 := "1";
    r3287 := "1";
    r3289 := (r3273 & r3275 & r3277 & r3279 & r3281 & r3283 & r3285 & r3287);
    r3291 := "1";
    r3293 := "1";
    r3295 := "0";
    r3297 := "1";
    r3299 := "0";
    r3301 := "1";
    r3303 := "1";
    r3305 := "1";
    r3307 := (r3291 & r3293 & r3295 & r3297 & r3299 & r3301 & r3303 & r3305);
    r3309 := "0";
    r3311 := "1";
    r3313 := "0";
    r3315 := "1";
    r3317 := "0";
    r3319 := "1";
    r3321 := "1";
    r3323 := "1";
    r3325 := (r3309 & r3311 & r3313 & r3315 & r3317 & r3319 & r3321 & r3323);
    r3327 := "1";
    r3329 := "0";
    r3331 := "0";
    r3333 := "1";
    r3335 := "0";
    r3337 := "1";
    r3339 := "1";
    r3341 := "1";
    r3343 := (r3327 & r3329 & r3331 & r3333 & r3335 & r3337 & r3339 & r3341);
    r3345 := "0";
    r3347 := "0";
    r3349 := "0";
    r3351 := "1";
    r3353 := "0";
    r3355 := "1";
    r3357 := "1";
    r3359 := "1";
    r3361 := (r3345 & r3347 & r3349 & r3351 & r3353 & r3355 & r3357 & r3359);
    r3363 := "1";
    r3365 := "1";
    r3367 := "1";
    r3369 := "0";
    r3371 := "0";
    r3373 := "1";
    r3375 := "1";
    r3377 := "1";
    r3379 := (r3363 & r3365 & r3367 & r3369 & r3371 & r3373 & r3375 & r3377);
    r3381 := "0";
    r3383 := "1";
    r3385 := "1";
    r3387 := "0";
    r3389 := "0";
    r3391 := "1";
    r3393 := "1";
    r3395 := "1";
    r3397 := (r3381 & r3383 & r3385 & r3387 & r3389 & r3391 & r3393 & r3395);
    r3399 := "1";
    r3401 := "0";
    r3403 := "1";
    r3405 := "0";
    r3407 := "0";
    r3409 := "1";
    r3411 := "1";
    r3413 := "1";
    r3415 := (r3399 & r3401 & r3403 & r3405 & r3407 & r3409 & r3411 & r3413);
    r3417 := "0";
    r3419 := "0";
    r3421 := "1";
    r3423 := "0";
    r3425 := "0";
    r3427 := "1";
    r3429 := "1";
    r3431 := "1";
    r3433 := (r3417 & r3419 & r3421 & r3423 & r3425 & r3427 & r3429 & r3431);
    r3435 := "1";
    r3437 := "1";
    r3439 := "0";
    r3441 := "0";
    r3443 := "0";
    r3445 := "1";
    r3447 := "1";
    r3449 := "1";
    r3451 := (r3435 & r3437 & r3439 & r3441 & r3443 & r3445 & r3447 & r3449);
    r3453 := "0";
    r3455 := "1";
    r3457 := "0";
    r3459 := "0";
    r3461 := "0";
    r3463 := "1";
    r3465 := "1";
    r3467 := "1";
    r3469 := (r3453 & r3455 & r3457 & r3459 & r3461 & r3463 & r3465 & r3467);
    r3471 := "1";
    r3473 := "0";
    r3475 := "0";
    r3477 := "0";
    r3479 := "0";
    r3481 := "1";
    r3483 := "1";
    r3485 := "1";
    r3487 := (r3471 & r3473 & r3475 & r3477 & r3479 & r3481 & r3483 & r3485);
    r3489 := "0";
    r3491 := "0";
    r3493 := "0";
    r3495 := "0";
    r3497 := "0";
    r3499 := "1";
    r3501 := "1";
    r3503 := "1";
    r3505 := (r3489 & r3491 & r3493 & r3495 & r3497 & r3499 & r3501 & r3503);
    r3507 := "1";
    r3509 := "1";
    r3511 := "1";
    r3513 := "1";
    r3515 := "1";
    r3517 := "0";
    r3519 := "1";
    r3521 := "1";
    r3523 := (r3507 & r3509 & r3511 & r3513 & r3515 & r3517 & r3519 & r3521);
    r3524 := (r3253 & r3271 & r3289 & r3307 & r3325 & r3343 & r3361 & r3379 & r3397 & r3415 & r3433 & r3451 & r3469 & r3487 & r3505 & r3523);
    return r3524;
  end rewire_key2_3233;
  function rewire_key1_2939 return std_logic_vector
  is
    variable r3230 : std_logic_vector(0 to 127) := (others => '0');
    variable r3229 : std_logic_vector(0 to 7) := (others => '0');
    variable r3227 : std_logic_vector(0 to 0) := (others => '0');
    variable r3225 : std_logic_vector(0 to 0) := (others => '0');
    variable r3223 : std_logic_vector(0 to 0) := (others => '0');
    variable r3221 : std_logic_vector(0 to 0) := (others => '0');
    variable r3219 : std_logic_vector(0 to 0) := (others => '0');
    variable r3217 : std_logic_vector(0 to 0) := (others => '0');
    variable r3215 : std_logic_vector(0 to 0) := (others => '0');
    variable r3213 : std_logic_vector(0 to 0) := (others => '0');
    variable r3211 : std_logic_vector(0 to 7) := (others => '0');
    variable r3209 : std_logic_vector(0 to 0) := (others => '0');
    variable r3207 : std_logic_vector(0 to 0) := (others => '0');
    variable r3205 : std_logic_vector(0 to 0) := (others => '0');
    variable r3203 : std_logic_vector(0 to 0) := (others => '0');
    variable r3201 : std_logic_vector(0 to 0) := (others => '0');
    variable r3199 : std_logic_vector(0 to 0) := (others => '0');
    variable r3197 : std_logic_vector(0 to 0) := (others => '0');
    variable r3195 : std_logic_vector(0 to 0) := (others => '0');
    variable r3193 : std_logic_vector(0 to 7) := (others => '0');
    variable r3191 : std_logic_vector(0 to 0) := (others => '0');
    variable r3189 : std_logic_vector(0 to 0) := (others => '0');
    variable r3187 : std_logic_vector(0 to 0) := (others => '0');
    variable r3185 : std_logic_vector(0 to 0) := (others => '0');
    variable r3183 : std_logic_vector(0 to 0) := (others => '0');
    variable r3181 : std_logic_vector(0 to 0) := (others => '0');
    variable r3179 : std_logic_vector(0 to 0) := (others => '0');
    variable r3177 : std_logic_vector(0 to 0) := (others => '0');
    variable r3175 : std_logic_vector(0 to 7) := (others => '0');
    variable r3173 : std_logic_vector(0 to 0) := (others => '0');
    variable r3171 : std_logic_vector(0 to 0) := (others => '0');
    variable r3169 : std_logic_vector(0 to 0) := (others => '0');
    variable r3167 : std_logic_vector(0 to 0) := (others => '0');
    variable r3165 : std_logic_vector(0 to 0) := (others => '0');
    variable r3163 : std_logic_vector(0 to 0) := (others => '0');
    variable r3161 : std_logic_vector(0 to 0) := (others => '0');
    variable r3159 : std_logic_vector(0 to 0) := (others => '0');
    variable r3157 : std_logic_vector(0 to 7) := (others => '0');
    variable r3155 : std_logic_vector(0 to 0) := (others => '0');
    variable r3153 : std_logic_vector(0 to 0) := (others => '0');
    variable r3151 : std_logic_vector(0 to 0) := (others => '0');
    variable r3149 : std_logic_vector(0 to 0) := (others => '0');
    variable r3147 : std_logic_vector(0 to 0) := (others => '0');
    variable r3145 : std_logic_vector(0 to 0) := (others => '0');
    variable r3143 : std_logic_vector(0 to 0) := (others => '0');
    variable r3141 : std_logic_vector(0 to 0) := (others => '0');
    variable r3139 : std_logic_vector(0 to 7) := (others => '0');
    variable r3137 : std_logic_vector(0 to 0) := (others => '0');
    variable r3135 : std_logic_vector(0 to 0) := (others => '0');
    variable r3133 : std_logic_vector(0 to 0) := (others => '0');
    variable r3131 : std_logic_vector(0 to 0) := (others => '0');
    variable r3129 : std_logic_vector(0 to 0) := (others => '0');
    variable r3127 : std_logic_vector(0 to 0) := (others => '0');
    variable r3125 : std_logic_vector(0 to 0) := (others => '0');
    variable r3123 : std_logic_vector(0 to 0) := (others => '0');
    variable r3121 : std_logic_vector(0 to 7) := (others => '0');
    variable r3119 : std_logic_vector(0 to 0) := (others => '0');
    variable r3117 : std_logic_vector(0 to 0) := (others => '0');
    variable r3115 : std_logic_vector(0 to 0) := (others => '0');
    variable r3113 : std_logic_vector(0 to 0) := (others => '0');
    variable r3111 : std_logic_vector(0 to 0) := (others => '0');
    variable r3109 : std_logic_vector(0 to 0) := (others => '0');
    variable r3107 : std_logic_vector(0 to 0) := (others => '0');
    variable r3105 : std_logic_vector(0 to 0) := (others => '0');
    variable r3103 : std_logic_vector(0 to 7) := (others => '0');
    variable r3101 : std_logic_vector(0 to 0) := (others => '0');
    variable r3099 : std_logic_vector(0 to 0) := (others => '0');
    variable r3097 : std_logic_vector(0 to 0) := (others => '0');
    variable r3095 : std_logic_vector(0 to 0) := (others => '0');
    variable r3093 : std_logic_vector(0 to 0) := (others => '0');
    variable r3091 : std_logic_vector(0 to 0) := (others => '0');
    variable r3089 : std_logic_vector(0 to 0) := (others => '0');
    variable r3087 : std_logic_vector(0 to 0) := (others => '0');
    variable r3085 : std_logic_vector(0 to 7) := (others => '0');
    variable r3083 : std_logic_vector(0 to 0) := (others => '0');
    variable r3081 : std_logic_vector(0 to 0) := (others => '0');
    variable r3079 : std_logic_vector(0 to 0) := (others => '0');
    variable r3077 : std_logic_vector(0 to 0) := (others => '0');
    variable r3075 : std_logic_vector(0 to 0) := (others => '0');
    variable r3073 : std_logic_vector(0 to 0) := (others => '0');
    variable r3071 : std_logic_vector(0 to 0) := (others => '0');
    variable r3069 : std_logic_vector(0 to 0) := (others => '0');
    variable r3067 : std_logic_vector(0 to 7) := (others => '0');
    variable r3065 : std_logic_vector(0 to 0) := (others => '0');
    variable r3063 : std_logic_vector(0 to 0) := (others => '0');
    variable r3061 : std_logic_vector(0 to 0) := (others => '0');
    variable r3059 : std_logic_vector(0 to 0) := (others => '0');
    variable r3057 : std_logic_vector(0 to 0) := (others => '0');
    variable r3055 : std_logic_vector(0 to 0) := (others => '0');
    variable r3053 : std_logic_vector(0 to 0) := (others => '0');
    variable r3051 : std_logic_vector(0 to 0) := (others => '0');
    variable r3049 : std_logic_vector(0 to 7) := (others => '0');
    variable r3047 : std_logic_vector(0 to 0) := (others => '0');
    variable r3045 : std_logic_vector(0 to 0) := (others => '0');
    variable r3043 : std_logic_vector(0 to 0) := (others => '0');
    variable r3041 : std_logic_vector(0 to 0) := (others => '0');
    variable r3039 : std_logic_vector(0 to 0) := (others => '0');
    variable r3037 : std_logic_vector(0 to 0) := (others => '0');
    variable r3035 : std_logic_vector(0 to 0) := (others => '0');
    variable r3033 : std_logic_vector(0 to 0) := (others => '0');
    variable r3031 : std_logic_vector(0 to 7) := (others => '0');
    variable r3029 : std_logic_vector(0 to 0) := (others => '0');
    variable r3027 : std_logic_vector(0 to 0) := (others => '0');
    variable r3025 : std_logic_vector(0 to 0) := (others => '0');
    variable r3023 : std_logic_vector(0 to 0) := (others => '0');
    variable r3021 : std_logic_vector(0 to 0) := (others => '0');
    variable r3019 : std_logic_vector(0 to 0) := (others => '0');
    variable r3017 : std_logic_vector(0 to 0) := (others => '0');
    variable r3015 : std_logic_vector(0 to 0) := (others => '0');
    variable r3013 : std_logic_vector(0 to 7) := (others => '0');
    variable r3011 : std_logic_vector(0 to 0) := (others => '0');
    variable r3009 : std_logic_vector(0 to 0) := (others => '0');
    variable r3007 : std_logic_vector(0 to 0) := (others => '0');
    variable r3005 : std_logic_vector(0 to 0) := (others => '0');
    variable r3003 : std_logic_vector(0 to 0) := (others => '0');
    variable r3001 : std_logic_vector(0 to 0) := (others => '0');
    variable r2999 : std_logic_vector(0 to 0) := (others => '0');
    variable r2997 : std_logic_vector(0 to 0) := (others => '0');
    variable r2995 : std_logic_vector(0 to 7) := (others => '0');
    variable r2993 : std_logic_vector(0 to 0) := (others => '0');
    variable r2991 : std_logic_vector(0 to 0) := (others => '0');
    variable r2989 : std_logic_vector(0 to 0) := (others => '0');
    variable r2987 : std_logic_vector(0 to 0) := (others => '0');
    variable r2985 : std_logic_vector(0 to 0) := (others => '0');
    variable r2983 : std_logic_vector(0 to 0) := (others => '0');
    variable r2981 : std_logic_vector(0 to 0) := (others => '0');
    variable r2979 : std_logic_vector(0 to 0) := (others => '0');
    variable r2977 : std_logic_vector(0 to 7) := (others => '0');
    variable r2975 : std_logic_vector(0 to 0) := (others => '0');
    variable r2973 : std_logic_vector(0 to 0) := (others => '0');
    variable r2971 : std_logic_vector(0 to 0) := (others => '0');
    variable r2969 : std_logic_vector(0 to 0) := (others => '0');
    variable r2967 : std_logic_vector(0 to 0) := (others => '0');
    variable r2965 : std_logic_vector(0 to 0) := (others => '0');
    variable r2963 : std_logic_vector(0 to 0) := (others => '0');
    variable r2961 : std_logic_vector(0 to 0) := (others => '0');
    variable r2959 : std_logic_vector(0 to 7) := (others => '0');
    variable r2957 : std_logic_vector(0 to 0) := (others => '0');
    variable r2955 : std_logic_vector(0 to 0) := (others => '0');
    variable r2953 : std_logic_vector(0 to 0) := (others => '0');
    variable r2951 : std_logic_vector(0 to 0) := (others => '0');
    variable r2949 : std_logic_vector(0 to 0) := (others => '0');
    variable r2947 : std_logic_vector(0 to 0) := (others => '0');
    variable r2945 : std_logic_vector(0 to 0) := (others => '0');
    variable r2943 : std_logic_vector(0 to 0) := (others => '0');
  begin
    r2943 := "0";
    r2945 := "1";
    r2947 := "1";
    r2949 := "1";
    r2951 := "1";
    r2953 := "1";
    r2955 := "1";
    r2957 := "1";
    r2959 := (r2943 & r2945 & r2947 & r2949 & r2951 & r2953 & r2955 & r2957);
    r2961 := "1";
    r2963 := "0";
    r2965 := "1";
    r2967 := "1";
    r2969 := "1";
    r2971 := "1";
    r2973 := "1";
    r2975 := "1";
    r2977 := (r2961 & r2963 & r2965 & r2967 & r2969 & r2971 & r2973 & r2975);
    r2979 := "0";
    r2981 := "0";
    r2983 := "1";
    r2985 := "1";
    r2987 := "1";
    r2989 := "1";
    r2991 := "1";
    r2993 := "1";
    r2995 := (r2979 & r2981 & r2983 & r2985 & r2987 & r2989 & r2991 & r2993);
    r2997 := "1";
    r2999 := "1";
    r3001 := "0";
    r3003 := "1";
    r3005 := "1";
    r3007 := "1";
    r3009 := "1";
    r3011 := "1";
    r3013 := (r2997 & r2999 & r3001 & r3003 & r3005 & r3007 & r3009 & r3011);
    r3015 := "0";
    r3017 := "1";
    r3019 := "0";
    r3021 := "1";
    r3023 := "1";
    r3025 := "1";
    r3027 := "1";
    r3029 := "1";
    r3031 := (r3015 & r3017 & r3019 & r3021 & r3023 & r3025 & r3027 & r3029);
    r3033 := "1";
    r3035 := "0";
    r3037 := "0";
    r3039 := "1";
    r3041 := "1";
    r3043 := "1";
    r3045 := "1";
    r3047 := "1";
    r3049 := (r3033 & r3035 & r3037 & r3039 & r3041 & r3043 & r3045 & r3047);
    r3051 := "0";
    r3053 := "0";
    r3055 := "0";
    r3057 := "1";
    r3059 := "1";
    r3061 := "1";
    r3063 := "1";
    r3065 := "1";
    r3067 := (r3051 & r3053 & r3055 & r3057 & r3059 & r3061 & r3063 & r3065);
    r3069 := "1";
    r3071 := "1";
    r3073 := "1";
    r3075 := "0";
    r3077 := "1";
    r3079 := "1";
    r3081 := "1";
    r3083 := "1";
    r3085 := (r3069 & r3071 & r3073 & r3075 & r3077 & r3079 & r3081 & r3083);
    r3087 := "0";
    r3089 := "1";
    r3091 := "1";
    r3093 := "0";
    r3095 := "1";
    r3097 := "1";
    r3099 := "1";
    r3101 := "1";
    r3103 := (r3087 & r3089 & r3091 & r3093 & r3095 & r3097 & r3099 & r3101);
    r3105 := "1";
    r3107 := "0";
    r3109 := "1";
    r3111 := "0";
    r3113 := "1";
    r3115 := "1";
    r3117 := "1";
    r3119 := "1";
    r3121 := (r3105 & r3107 & r3109 & r3111 & r3113 & r3115 & r3117 & r3119);
    r3123 := "0";
    r3125 := "0";
    r3127 := "1";
    r3129 := "0";
    r3131 := "1";
    r3133 := "1";
    r3135 := "1";
    r3137 := "1";
    r3139 := (r3123 & r3125 & r3127 & r3129 & r3131 & r3133 & r3135 & r3137);
    r3141 := "1";
    r3143 := "1";
    r3145 := "0";
    r3147 := "0";
    r3149 := "1";
    r3151 := "1";
    r3153 := "1";
    r3155 := "1";
    r3157 := (r3141 & r3143 & r3145 & r3147 & r3149 & r3151 & r3153 & r3155);
    r3159 := "0";
    r3161 := "1";
    r3163 := "0";
    r3165 := "0";
    r3167 := "1";
    r3169 := "1";
    r3171 := "1";
    r3173 := "1";
    r3175 := (r3159 & r3161 & r3163 & r3165 & r3167 & r3169 & r3171 & r3173);
    r3177 := "1";
    r3179 := "0";
    r3181 := "0";
    r3183 := "0";
    r3185 := "1";
    r3187 := "1";
    r3189 := "1";
    r3191 := "1";
    r3193 := (r3177 & r3179 & r3181 & r3183 & r3185 & r3187 & r3189 & r3191);
    r3195 := "0";
    r3197 := "0";
    r3199 := "0";
    r3201 := "0";
    r3203 := "1";
    r3205 := "1";
    r3207 := "1";
    r3209 := "1";
    r3211 := (r3195 & r3197 & r3199 & r3201 & r3203 & r3205 & r3207 & r3209);
    r3213 := "1";
    r3215 := "1";
    r3217 := "1";
    r3219 := "1";
    r3221 := "0";
    r3223 := "1";
    r3225 := "1";
    r3227 := "1";
    r3229 := (r3213 & r3215 & r3217 & r3219 & r3221 & r3223 & r3225 & r3227);
    r3230 := (r2959 & r2977 & r2995 & r3013 & r3031 & r3049 & r3067 & r3085 & r3103 & r3121 & r3139 & r3157 & r3175 & r3193 & r3211 & r3229);
    return r3230;
  end rewire_key1_2939;
  function rewire_buildSalsa256_1182(r1183 : std_logic_vector ; r1184 : std_logic_vector ; r1185 : std_logic_vector ; r1186 : std_logic_vector) return std_logic_vector
  is
    variable r2938 : std_logic_vector(0 to 511) := (others => '0');
    variable r2937 : std_logic_vector(0 to 511) := (others => '0');
    variable r1660 : std_logic_vector(0 to 511) := (others => '0');
    variable r1659 : std_logic_vector(0 to 511) := (others => '0');
    variable b1657 : boolean := false;
    variable b1656 : boolean := false;
    variable b1655 : boolean := false;
    variable b1654 : boolean := false;
    variable b1653 : boolean := false;
    variable b1652 : boolean := false;
    variable r1651 : std_logic_vector(0 to 7) := (others => '0');
    variable r1650 : std_logic_vector(0 to 7) := (others => '0');
    variable r1649 : std_logic_vector(0 to 7) := (others => '0');
    variable r1648 : std_logic_vector(0 to 7) := (others => '0');
    variable b1647 : boolean := false;
    variable b1646 : boolean := false;
    variable b1645 : boolean := false;
    variable b1644 : boolean := false;
    variable b1643 : boolean := false;
    variable b1642 : boolean := false;
    variable r1641 : std_logic_vector(0 to 7) := (others => '0');
    variable r1640 : std_logic_vector(0 to 7) := (others => '0');
    variable r1639 : std_logic_vector(0 to 7) := (others => '0');
    variable r1638 : std_logic_vector(0 to 7) := (others => '0');
    variable b1637 : boolean := false;
    variable b1636 : boolean := false;
    variable b1635 : boolean := false;
    variable b1634 : boolean := false;
    variable b1633 : boolean := false;
    variable b1632 : boolean := false;
    variable r1631 : std_logic_vector(0 to 7) := (others => '0');
    variable r1630 : std_logic_vector(0 to 7) := (others => '0');
    variable r1629 : std_logic_vector(0 to 7) := (others => '0');
    variable r1628 : std_logic_vector(0 to 7) := (others => '0');
    variable b1627 : boolean := false;
    variable b1626 : boolean := false;
    variable b1625 : boolean := false;
    variable b1624 : boolean := false;
    variable b1623 : boolean := false;
    variable b1622 : boolean := false;
    variable r1621 : std_logic_vector(0 to 7) := (others => '0');
    variable r1620 : std_logic_vector(0 to 7) := (others => '0');
    variable r1619 : std_logic_vector(0 to 7) := (others => '0');
    variable r1618 : std_logic_vector(0 to 7) := (others => '0');
    variable b1617 : boolean := false;
    variable r1616 : std_logic_vector(0 to 31) := (others => '0');
    variable r1615 : std_logic_vector(0 to 31) := (others => '0');
    variable r1614 : std_logic_vector(0 to 31) := (others => '0');
    variable r1613 : std_logic_vector(0 to 31) := (others => '0');
    variable b1612 : boolean := false;
    variable r1611 : std_logic_vector(0 to 511) := (others => '0');
    variable r1610 : std_logic_vector(0 to 127) := (others => '0');
    variable r1609 : std_logic_vector(0 to 31) := (others => '0');
    variable r1534 : std_logic_vector(0 to 31) := (others => '0');
    variable r1532 : std_logic_vector(0 to 31) := (others => '0');
    variable r1457 : std_logic_vector(0 to 31) := (others => '0');
    variable r1455 : std_logic_vector(0 to 31) := (others => '0');
    variable r1380 : std_logic_vector(0 to 31) := (others => '0');
    variable r1378 : std_logic_vector(0 to 31) := (others => '0');
    variable r1303 : std_logic_vector(0 to 31) := (others => '0');
    variable b1300 : boolean := false;
    variable b1299 : boolean := false;
    variable b1298 : boolean := false;
    variable b1297 : boolean := false;
    variable b1296 : boolean := false;
    variable b1295 : boolean := false;
    variable b1294 : boolean := false;
    variable b1293 : boolean := false;
    variable b1292 : boolean := false;
    variable b1291 : boolean := false;
    variable r1290 : std_logic_vector(0 to 7) := (others => '0');
    variable r1289 : std_logic_vector(0 to 7) := (others => '0');
    variable r1288 : std_logic_vector(0 to 7) := (others => '0');
    variable r1287 : std_logic_vector(0 to 7) := (others => '0');
    variable r1286 : std_logic_vector(0 to 7) := (others => '0');
    variable r1285 : std_logic_vector(0 to 7) := (others => '0');
    variable r1284 : std_logic_vector(0 to 7) := (others => '0');
    variable r1283 : std_logic_vector(0 to 7) := (others => '0');
    variable b1282 : boolean := false;
    variable b1281 : boolean := false;
    variable b1280 : boolean := false;
    variable b1279 : boolean := false;
    variable b1278 : boolean := false;
    variable b1277 : boolean := false;
    variable b1276 : boolean := false;
    variable b1275 : boolean := false;
    variable b1274 : boolean := false;
    variable b1273 : boolean := false;
    variable r1272 : std_logic_vector(0 to 7) := (others => '0');
    variable r1271 : std_logic_vector(0 to 7) := (others => '0');
    variable r1270 : std_logic_vector(0 to 7) := (others => '0');
    variable r1269 : std_logic_vector(0 to 7) := (others => '0');
    variable r1268 : std_logic_vector(0 to 7) := (others => '0');
    variable r1267 : std_logic_vector(0 to 7) := (others => '0');
    variable r1266 : std_logic_vector(0 to 7) := (others => '0');
    variable r1265 : std_logic_vector(0 to 7) := (others => '0');
    variable b1264 : boolean := false;
    variable b1263 : boolean := false;
    variable b1262 : boolean := false;
    variable b1261 : boolean := false;
    variable b1260 : boolean := false;
    variable b1259 : boolean := false;
    variable b1258 : boolean := false;
    variable b1257 : boolean := false;
    variable b1256 : boolean := false;
    variable b1255 : boolean := false;
    variable b1254 : boolean := false;
    variable b1253 : boolean := false;
    variable b1252 : boolean := false;
    variable b1251 : boolean := false;
    variable b1250 : boolean := false;
    variable b1249 : boolean := false;
    variable b1248 : boolean := false;
    variable b1247 : boolean := false;
    variable r1246 : std_logic_vector(0 to 7) := (others => '0');
    variable r1245 : std_logic_vector(0 to 7) := (others => '0');
    variable r1244 : std_logic_vector(0 to 7) := (others => '0');
    variable r1243 : std_logic_vector(0 to 7) := (others => '0');
    variable r1242 : std_logic_vector(0 to 7) := (others => '0');
    variable r1241 : std_logic_vector(0 to 7) := (others => '0');
    variable r1240 : std_logic_vector(0 to 7) := (others => '0');
    variable r1239 : std_logic_vector(0 to 7) := (others => '0');
    variable r1238 : std_logic_vector(0 to 7) := (others => '0');
    variable r1237 : std_logic_vector(0 to 7) := (others => '0');
    variable r1236 : std_logic_vector(0 to 7) := (others => '0');
    variable r1235 : std_logic_vector(0 to 7) := (others => '0');
    variable r1234 : std_logic_vector(0 to 7) := (others => '0');
    variable r1233 : std_logic_vector(0 to 7) := (others => '0');
    variable r1232 : std_logic_vector(0 to 7) := (others => '0');
    variable r1231 : std_logic_vector(0 to 7) := (others => '0');
    variable b1230 : boolean := false;
    variable b1229 : boolean := false;
    variable b1228 : boolean := false;
    variable b1227 : boolean := false;
    variable b1226 : boolean := false;
    variable b1225 : boolean := false;
    variable b1224 : boolean := false;
    variable b1223 : boolean := false;
    variable b1222 : boolean := false;
    variable b1221 : boolean := false;
    variable b1220 : boolean := false;
    variable b1219 : boolean := false;
    variable b1218 : boolean := false;
    variable b1217 : boolean := false;
    variable b1216 : boolean := false;
    variable b1215 : boolean := false;
    variable b1214 : boolean := false;
    variable b1213 : boolean := false;
    variable r1212 : std_logic_vector(0 to 7) := (others => '0');
    variable r1211 : std_logic_vector(0 to 7) := (others => '0');
    variable r1210 : std_logic_vector(0 to 7) := (others => '0');
    variable r1209 : std_logic_vector(0 to 7) := (others => '0');
    variable r1208 : std_logic_vector(0 to 7) := (others => '0');
    variable r1207 : std_logic_vector(0 to 7) := (others => '0');
    variable r1206 : std_logic_vector(0 to 7) := (others => '0');
    variable r1205 : std_logic_vector(0 to 7) := (others => '0');
    variable r1204 : std_logic_vector(0 to 7) := (others => '0');
    variable r1203 : std_logic_vector(0 to 7) := (others => '0');
    variable r1202 : std_logic_vector(0 to 7) := (others => '0');
    variable r1201 : std_logic_vector(0 to 7) := (others => '0');
    variable r1200 : std_logic_vector(0 to 7) := (others => '0');
    variable r1199 : std_logic_vector(0 to 7) := (others => '0');
    variable r1198 : std_logic_vector(0 to 7) := (others => '0');
    variable r1197 : std_logic_vector(0 to 7) := (others => '0');
    variable b1196 : boolean := false;
    variable r1195 : std_logic_vector(0 to 63) := (others => '0');
    variable r1194 : std_logic_vector(0 to 63) := (others => '0');
    variable r1193 : std_logic_vector(0 to 127) := (others => '0');
    variable r1192 : std_logic_vector(0 to 127) := (others => '0');
    variable b1191 : boolean := false;
    variable r1190 : std_logic_vector(0 to 511) := (others => '0');
    variable r1189 : std_logic_vector(0 to 383) := (others => '0');
  begin
    b1191 := true;
    r1192 := r1189(0 to 127);
    r1193 := r1189(128 to 255);
    r1194 := r1189(256 to 319);
    r1195 := r1189(320 to 383);
    b1196 := true;
    r1197 := r1192(0 to 7);
    r1198 := r1192(8 to 15);
    r1199 := r1192(16 to 23);
    r1200 := r1192(24 to 31);
    r1201 := r1192(32 to 39);
    r1202 := r1192(40 to 47);
    r1203 := r1192(48 to 55);
    r1204 := r1192(56 to 63);
    r1205 := r1192(64 to 71);
    r1206 := r1192(72 to 79);
    r1207 := r1192(80 to 87);
    r1208 := r1192(88 to 95);
    r1209 := r1192(96 to 103);
    r1210 := r1192(104 to 111);
    r1211 := r1192(112 to 119);
    r1212 := r1192(120 to 127);
    b1213 := true;
    b1214 := true;
    b1215 := true;
    b1216 := true;
    b1217 := true;
    b1218 := true;
    b1219 := true;
    b1220 := true;
    b1221 := true;
    b1222 := true;
    b1223 := true;
    b1224 := true;
    b1225 := true;
    b1226 := true;
    b1227 := true;
    b1228 := true;
    b1229 := (b1213 AND (b1214 AND (b1215 AND (b1216 AND (b1217 AND (b1218 AND (b1219 AND (b1220 AND (b1221 AND (b1222 AND (b1223 AND (b1224 AND (b1225 AND (b1226 AND (b1227 AND b1228)))))))))))))));
    b1230 := true;
    r1231 := r1193(0 to 7);
    r1232 := r1193(8 to 15);
    r1233 := r1193(16 to 23);
    r1234 := r1193(24 to 31);
    r1235 := r1193(32 to 39);
    r1236 := r1193(40 to 47);
    r1237 := r1193(48 to 55);
    r1238 := r1193(56 to 63);
    r1239 := r1193(64 to 71);
    r1240 := r1193(72 to 79);
    r1241 := r1193(80 to 87);
    r1242 := r1193(88 to 95);
    r1243 := r1193(96 to 103);
    r1244 := r1193(104 to 111);
    r1245 := r1193(112 to 119);
    r1246 := r1193(120 to 127);
    b1247 := true;
    b1248 := true;
    b1249 := true;
    b1250 := true;
    b1251 := true;
    b1252 := true;
    b1253 := true;
    b1254 := true;
    b1255 := true;
    b1256 := true;
    b1257 := true;
    b1258 := true;
    b1259 := true;
    b1260 := true;
    b1261 := true;
    b1262 := true;
    b1263 := (b1247 AND (b1248 AND (b1249 AND (b1250 AND (b1251 AND (b1252 AND (b1253 AND (b1254 AND (b1255 AND (b1256 AND (b1257 AND (b1258 AND (b1259 AND (b1260 AND (b1261 AND b1262)))))))))))))));
    b1264 := true;
    r1265 := r1194(0 to 7);
    r1266 := r1194(8 to 15);
    r1267 := r1194(16 to 23);
    r1268 := r1194(24 to 31);
    r1269 := r1194(32 to 39);
    r1270 := r1194(40 to 47);
    r1271 := r1194(48 to 55);
    r1272 := r1194(56 to 63);
    b1273 := true;
    b1274 := true;
    b1275 := true;
    b1276 := true;
    b1277 := true;
    b1278 := true;
    b1279 := true;
    b1280 := true;
    b1281 := (b1273 AND (b1274 AND (b1275 AND (b1276 AND (b1277 AND (b1278 AND (b1279 AND b1280)))))));
    b1282 := true;
    r1283 := r1195(0 to 7);
    r1284 := r1195(8 to 15);
    r1285 := r1195(16 to 23);
    r1286 := r1195(24 to 31);
    r1287 := r1195(32 to 39);
    r1288 := r1195(40 to 47);
    r1289 := r1195(48 to 55);
    r1290 := r1195(56 to 63);
    b1291 := true;
    b1292 := true;
    b1293 := true;
    b1294 := true;
    b1295 := true;
    b1296 := true;
    b1297 := true;
    b1298 := true;
    b1299 := (b1291 AND (b1292 AND (b1293 AND (b1294 AND (b1295 AND (b1296 AND (b1297 AND b1298)))))));
    b1300 := (b1229 AND (b1263 AND (b1281 AND b1299)));
    if b1300 then
      b1612 := true;
      r1613 := r1610(0 to 31);
      r1614 := r1610(32 to 63);
      r1615 := r1610(64 to 95);
      r1616 := r1610(96 to 127);
      b1617 := true;
      r1618 := r1613(0 to 7);
      r1619 := r1613(8 to 15);
      r1620 := r1613(16 to 23);
      r1621 := r1613(24 to 31);
      b1622 := true;
      b1623 := true;
      b1624 := true;
      b1625 := true;
      b1626 := (b1622 AND (b1623 AND (b1624 AND b1625)));
      b1627 := true;
      r1628 := r1614(0 to 7);
      r1629 := r1614(8 to 15);
      r1630 := r1614(16 to 23);
      r1631 := r1614(24 to 31);
      b1632 := true;
      b1633 := true;
      b1634 := true;
      b1635 := true;
      b1636 := (b1632 AND (b1633 AND (b1634 AND b1635)));
      b1637 := true;
      r1638 := r1615(0 to 7);
      r1639 := r1615(8 to 15);
      r1640 := r1615(16 to 23);
      r1641 := r1615(24 to 31);
      b1642 := true;
      b1643 := true;
      b1644 := true;
      b1645 := true;
      b1646 := (b1642 AND (b1643 AND (b1644 AND b1645)));
      b1647 := true;
      r1648 := r1616(0 to 7);
      r1649 := r1616(8 to 15);
      r1650 := r1616(16 to 23);
      r1651 := r1616(24 to 31);
      b1652 := true;
      b1653 := true;
      b1654 := true;
      b1655 := true;
      b1656 := (b1652 AND (b1653 AND (b1654 AND b1655)));
      b1657 := (b1626 AND (b1636 AND (b1646 AND b1656)));
      if b1657 then
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        r2937 := (r1618 & r1619 & r1620 & r1621 & r1197 & r1198 & r1199 & r1200 & r1201 & r1202 & r1203 & r1204 & r1205 & r1206 & r1207 & r1208 & r1209 & r1210 & r1211 & r1212 & r1628 & r1629 & r1630 & r1631 & r1265 & r1266 & r1267 & r1268 & r1269 & r1270 & r1271 & r1272 & r1283 & r1284 & r1285 & r1286 & r1287 & r1288 & r1289 & r1290 & r1638 & r1639 & r1640 & r1641 & r1231 & r1232 & r1233 & r1234 & r1235 & r1236 & r1237 & r1238 & r1239 & r1240 & r1241 & r1242 & r1243 & r1244 & r1245 & r1246 & r1648 & r1649 & r1650 & r1651);
        r2938 := rewire_salsaHash_1658(r2937);
        r1611 := r2938;
      end if;
      r1190 := r1611;
    end if;
    return r1190;
  end rewire_buildSalsa256_1182;
  function rewire_salsaHash_1658(r1659 : std_logic_vector) return std_logic_vector
  is
    variable r2935 : std_logic_vector(0 to 511) := (others => '0');
    variable r2934 : std_logic_vector(0 to 511) := (others => '0');
    variable r2933 : std_logic_vector(0 to 511) := (others => '0');
    variable r2604 : std_logic_vector(0 to 511) := (others => '0');
    variable r2603 : std_logic_vector(0 to 511) := (others => '0');
    variable r1980 : std_logic_vector(0 to 511) := (others => '0');
    variable r1979 : std_logic_vector(0 to 511) := (others => '0');
    variable r1663 : std_logic_vector(0 to 511) := (others => '0');
    variable r1662 : std_logic_vector(0 to 511) := (others => '0');
  begin
    null;
    r2933 := rewire_impwords_2602(r1659);
    r2934 := rewire_salsaHashp_1978(r2933);
    r2935 := rewire_expwords_1661(r2934);
    return r2935;
  end rewire_salsaHash_1658;
  function rewire_impwords_2602(r2603 : std_logic_vector) return std_logic_vector
  is
    variable r2932 : std_logic_vector(0 to 511) := (others => '0');
    variable r2930 : std_logic_vector(0 to 31) := (others => '0');
    variable r2929 : std_logic_vector(0 to 31) := (others => '0');
    variable r2927 : std_logic_vector(0 to 31) := (others => '0');
    variable r2926 : std_logic_vector(0 to 31) := (others => '0');
    variable r2924 : std_logic_vector(0 to 31) := (others => '0');
    variable r2923 : std_logic_vector(0 to 31) := (others => '0');
    variable r2921 : std_logic_vector(0 to 31) := (others => '0');
    variable r2920 : std_logic_vector(0 to 31) := (others => '0');
    variable r2918 : std_logic_vector(0 to 31) := (others => '0');
    variable r2917 : std_logic_vector(0 to 31) := (others => '0');
    variable r2915 : std_logic_vector(0 to 31) := (others => '0');
    variable r2914 : std_logic_vector(0 to 31) := (others => '0');
    variable r2912 : std_logic_vector(0 to 31) := (others => '0');
    variable r2911 : std_logic_vector(0 to 31) := (others => '0');
    variable r2909 : std_logic_vector(0 to 31) := (others => '0');
    variable r2908 : std_logic_vector(0 to 31) := (others => '0');
    variable r2906 : std_logic_vector(0 to 31) := (others => '0');
    variable r2905 : std_logic_vector(0 to 31) := (others => '0');
    variable r2903 : std_logic_vector(0 to 31) := (others => '0');
    variable r2902 : std_logic_vector(0 to 31) := (others => '0');
    variable r2900 : std_logic_vector(0 to 31) := (others => '0');
    variable r2899 : std_logic_vector(0 to 31) := (others => '0');
    variable r2897 : std_logic_vector(0 to 31) := (others => '0');
    variable r2896 : std_logic_vector(0 to 31) := (others => '0');
    variable r2894 : std_logic_vector(0 to 31) := (others => '0');
    variable r2893 : std_logic_vector(0 to 31) := (others => '0');
    variable r2891 : std_logic_vector(0 to 31) := (others => '0');
    variable r2890 : std_logic_vector(0 to 31) := (others => '0');
    variable r2888 : std_logic_vector(0 to 31) := (others => '0');
    variable r2887 : std_logic_vector(0 to 31) := (others => '0');
    variable r2885 : std_logic_vector(0 to 31) := (others => '0');
    variable r2884 : std_logic_vector(0 to 31) := (others => '0');
    variable r2738 : std_logic_vector(0 to 31) := (others => '0');
    variable r2737 : std_logic_vector(0 to 31) := (others => '0');
    variable b2735 : boolean := false;
    variable b2734 : boolean := false;
    variable b2733 : boolean := false;
    variable b2732 : boolean := false;
    variable b2731 : boolean := false;
    variable b2730 : boolean := false;
    variable b2729 : boolean := false;
    variable b2728 : boolean := false;
    variable b2727 : boolean := false;
    variable b2726 : boolean := false;
    variable b2725 : boolean := false;
    variable b2724 : boolean := false;
    variable b2723 : boolean := false;
    variable b2722 : boolean := false;
    variable b2721 : boolean := false;
    variable b2720 : boolean := false;
    variable b2719 : boolean := false;
    variable b2718 : boolean := false;
    variable b2717 : boolean := false;
    variable b2716 : boolean := false;
    variable b2715 : boolean := false;
    variable b2714 : boolean := false;
    variable b2713 : boolean := false;
    variable b2712 : boolean := false;
    variable b2711 : boolean := false;
    variable b2710 : boolean := false;
    variable b2709 : boolean := false;
    variable b2708 : boolean := false;
    variable b2707 : boolean := false;
    variable b2706 : boolean := false;
    variable b2705 : boolean := false;
    variable b2704 : boolean := false;
    variable b2703 : boolean := false;
    variable b2702 : boolean := false;
    variable b2701 : boolean := false;
    variable b2700 : boolean := false;
    variable b2699 : boolean := false;
    variable b2698 : boolean := false;
    variable b2697 : boolean := false;
    variable b2696 : boolean := false;
    variable b2695 : boolean := false;
    variable b2694 : boolean := false;
    variable b2693 : boolean := false;
    variable b2692 : boolean := false;
    variable b2691 : boolean := false;
    variable b2690 : boolean := false;
    variable b2689 : boolean := false;
    variable b2688 : boolean := false;
    variable b2687 : boolean := false;
    variable b2686 : boolean := false;
    variable b2685 : boolean := false;
    variable b2684 : boolean := false;
    variable b2683 : boolean := false;
    variable b2682 : boolean := false;
    variable b2681 : boolean := false;
    variable b2680 : boolean := false;
    variable b2679 : boolean := false;
    variable b2678 : boolean := false;
    variable b2677 : boolean := false;
    variable b2676 : boolean := false;
    variable b2675 : boolean := false;
    variable b2674 : boolean := false;
    variable b2673 : boolean := false;
    variable b2672 : boolean := false;
    variable b2671 : boolean := false;
    variable r2670 : std_logic_vector(0 to 7) := (others => '0');
    variable r2669 : std_logic_vector(0 to 7) := (others => '0');
    variable r2668 : std_logic_vector(0 to 7) := (others => '0');
    variable r2667 : std_logic_vector(0 to 7) := (others => '0');
    variable r2666 : std_logic_vector(0 to 7) := (others => '0');
    variable r2665 : std_logic_vector(0 to 7) := (others => '0');
    variable r2664 : std_logic_vector(0 to 7) := (others => '0');
    variable r2663 : std_logic_vector(0 to 7) := (others => '0');
    variable r2662 : std_logic_vector(0 to 7) := (others => '0');
    variable r2661 : std_logic_vector(0 to 7) := (others => '0');
    variable r2660 : std_logic_vector(0 to 7) := (others => '0');
    variable r2659 : std_logic_vector(0 to 7) := (others => '0');
    variable r2658 : std_logic_vector(0 to 7) := (others => '0');
    variable r2657 : std_logic_vector(0 to 7) := (others => '0');
    variable r2656 : std_logic_vector(0 to 7) := (others => '0');
    variable r2655 : std_logic_vector(0 to 7) := (others => '0');
    variable r2654 : std_logic_vector(0 to 7) := (others => '0');
    variable r2653 : std_logic_vector(0 to 7) := (others => '0');
    variable r2652 : std_logic_vector(0 to 7) := (others => '0');
    variable r2651 : std_logic_vector(0 to 7) := (others => '0');
    variable r2650 : std_logic_vector(0 to 7) := (others => '0');
    variable r2649 : std_logic_vector(0 to 7) := (others => '0');
    variable r2648 : std_logic_vector(0 to 7) := (others => '0');
    variable r2647 : std_logic_vector(0 to 7) := (others => '0');
    variable r2646 : std_logic_vector(0 to 7) := (others => '0');
    variable r2645 : std_logic_vector(0 to 7) := (others => '0');
    variable r2644 : std_logic_vector(0 to 7) := (others => '0');
    variable r2643 : std_logic_vector(0 to 7) := (others => '0');
    variable r2642 : std_logic_vector(0 to 7) := (others => '0');
    variable r2641 : std_logic_vector(0 to 7) := (others => '0');
    variable r2640 : std_logic_vector(0 to 7) := (others => '0');
    variable r2639 : std_logic_vector(0 to 7) := (others => '0');
    variable r2638 : std_logic_vector(0 to 7) := (others => '0');
    variable r2637 : std_logic_vector(0 to 7) := (others => '0');
    variable r2636 : std_logic_vector(0 to 7) := (others => '0');
    variable r2635 : std_logic_vector(0 to 7) := (others => '0');
    variable r2634 : std_logic_vector(0 to 7) := (others => '0');
    variable r2633 : std_logic_vector(0 to 7) := (others => '0');
    variable r2632 : std_logic_vector(0 to 7) := (others => '0');
    variable r2631 : std_logic_vector(0 to 7) := (others => '0');
    variable r2630 : std_logic_vector(0 to 7) := (others => '0');
    variable r2629 : std_logic_vector(0 to 7) := (others => '0');
    variable r2628 : std_logic_vector(0 to 7) := (others => '0');
    variable r2627 : std_logic_vector(0 to 7) := (others => '0');
    variable r2626 : std_logic_vector(0 to 7) := (others => '0');
    variable r2625 : std_logic_vector(0 to 7) := (others => '0');
    variable r2624 : std_logic_vector(0 to 7) := (others => '0');
    variable r2623 : std_logic_vector(0 to 7) := (others => '0');
    variable r2622 : std_logic_vector(0 to 7) := (others => '0');
    variable r2621 : std_logic_vector(0 to 7) := (others => '0');
    variable r2620 : std_logic_vector(0 to 7) := (others => '0');
    variable r2619 : std_logic_vector(0 to 7) := (others => '0');
    variable r2618 : std_logic_vector(0 to 7) := (others => '0');
    variable r2617 : std_logic_vector(0 to 7) := (others => '0');
    variable r2616 : std_logic_vector(0 to 7) := (others => '0');
    variable r2615 : std_logic_vector(0 to 7) := (others => '0');
    variable r2614 : std_logic_vector(0 to 7) := (others => '0');
    variable r2613 : std_logic_vector(0 to 7) := (others => '0');
    variable r2612 : std_logic_vector(0 to 7) := (others => '0');
    variable r2611 : std_logic_vector(0 to 7) := (others => '0');
    variable r2610 : std_logic_vector(0 to 7) := (others => '0');
    variable r2609 : std_logic_vector(0 to 7) := (others => '0');
    variable r2608 : std_logic_vector(0 to 7) := (others => '0');
    variable r2607 : std_logic_vector(0 to 7) := (others => '0');
    variable b2606 : boolean := false;
    variable r2605 : std_logic_vector(0 to 511) := (others => '0');
  begin
    b2606 := true;
    r2607 := r2603(0 to 7);
    r2608 := r2603(8 to 15);
    r2609 := r2603(16 to 23);
    r2610 := r2603(24 to 31);
    r2611 := r2603(32 to 39);
    r2612 := r2603(40 to 47);
    r2613 := r2603(48 to 55);
    r2614 := r2603(56 to 63);
    r2615 := r2603(64 to 71);
    r2616 := r2603(72 to 79);
    r2617 := r2603(80 to 87);
    r2618 := r2603(88 to 95);
    r2619 := r2603(96 to 103);
    r2620 := r2603(104 to 111);
    r2621 := r2603(112 to 119);
    r2622 := r2603(120 to 127);
    r2623 := r2603(128 to 135);
    r2624 := r2603(136 to 143);
    r2625 := r2603(144 to 151);
    r2626 := r2603(152 to 159);
    r2627 := r2603(160 to 167);
    r2628 := r2603(168 to 175);
    r2629 := r2603(176 to 183);
    r2630 := r2603(184 to 191);
    r2631 := r2603(192 to 199);
    r2632 := r2603(200 to 207);
    r2633 := r2603(208 to 215);
    r2634 := r2603(216 to 223);
    r2635 := r2603(224 to 231);
    r2636 := r2603(232 to 239);
    r2637 := r2603(240 to 247);
    r2638 := r2603(248 to 255);
    r2639 := r2603(256 to 263);
    r2640 := r2603(264 to 271);
    r2641 := r2603(272 to 279);
    r2642 := r2603(280 to 287);
    r2643 := r2603(288 to 295);
    r2644 := r2603(296 to 303);
    r2645 := r2603(304 to 311);
    r2646 := r2603(312 to 319);
    r2647 := r2603(320 to 327);
    r2648 := r2603(328 to 335);
    r2649 := r2603(336 to 343);
    r2650 := r2603(344 to 351);
    r2651 := r2603(352 to 359);
    r2652 := r2603(360 to 367);
    r2653 := r2603(368 to 375);
    r2654 := r2603(376 to 383);
    r2655 := r2603(384 to 391);
    r2656 := r2603(392 to 399);
    r2657 := r2603(400 to 407);
    r2658 := r2603(408 to 415);
    r2659 := r2603(416 to 423);
    r2660 := r2603(424 to 431);
    r2661 := r2603(432 to 439);
    r2662 := r2603(440 to 447);
    r2663 := r2603(448 to 455);
    r2664 := r2603(456 to 463);
    r2665 := r2603(464 to 471);
    r2666 := r2603(472 to 479);
    r2667 := r2603(480 to 487);
    r2668 := r2603(488 to 495);
    r2669 := r2603(496 to 503);
    r2670 := r2603(504 to 511);
    b2671 := true;
    b2672 := true;
    b2673 := true;
    b2674 := true;
    b2675 := true;
    b2676 := true;
    b2677 := true;
    b2678 := true;
    b2679 := true;
    b2680 := true;
    b2681 := true;
    b2682 := true;
    b2683 := true;
    b2684 := true;
    b2685 := true;
    b2686 := true;
    b2687 := true;
    b2688 := true;
    b2689 := true;
    b2690 := true;
    b2691 := true;
    b2692 := true;
    b2693 := true;
    b2694 := true;
    b2695 := true;
    b2696 := true;
    b2697 := true;
    b2698 := true;
    b2699 := true;
    b2700 := true;
    b2701 := true;
    b2702 := true;
    b2703 := true;
    b2704 := true;
    b2705 := true;
    b2706 := true;
    b2707 := true;
    b2708 := true;
    b2709 := true;
    b2710 := true;
    b2711 := true;
    b2712 := true;
    b2713 := true;
    b2714 := true;
    b2715 := true;
    b2716 := true;
    b2717 := true;
    b2718 := true;
    b2719 := true;
    b2720 := true;
    b2721 := true;
    b2722 := true;
    b2723 := true;
    b2724 := true;
    b2725 := true;
    b2726 := true;
    b2727 := true;
    b2728 := true;
    b2729 := true;
    b2730 := true;
    b2731 := true;
    b2732 := true;
    b2733 := true;
    b2734 := true;
    b2735 := (b2671 AND (b2672 AND (b2673 AND (b2674 AND (b2675 AND (b2676 AND (b2677 AND (b2678 AND (b2679 AND (b2680 AND (b2681 AND (b2682 AND (b2683 AND (b2684 AND (b2685 AND (b2686 AND (b2687 AND (b2688 AND (b2689 AND (b2690 AND (b2691 AND (b2692 AND (b2693 AND (b2694 AND (b2695 AND (b2696 AND (b2697 AND (b2698 AND (b2699 AND (b2700 AND (b2701 AND (b2702 AND (b2703 AND (b2704 AND (b2705 AND (b2706 AND (b2707 AND (b2708 AND (b2709 AND (b2710 AND (b2711 AND (b2712 AND (b2713 AND (b2714 AND (b2715 AND (b2716 AND (b2717 AND (b2718 AND (b2719 AND (b2720 AND (b2721 AND (b2722 AND (b2723 AND (b2724 AND (b2725 AND (b2726 AND (b2727 AND (b2728 AND (b2729 AND (b2730 AND (b2731 AND (b2732 AND (b2733 AND b2734)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
    if b2735 then
      null;
      null;
      null;
      null;
      r2884 := (r2607 & r2608 & r2609 & r2610);
      r2885 := rewire_littleendian_2736(r2884);
      null;
      null;
      null;
      null;
      r2887 := (r2611 & r2612 & r2613 & r2614);
      r2888 := rewire_littleendian_2736(r2887);
      null;
      null;
      null;
      null;
      r2890 := (r2615 & r2616 & r2617 & r2618);
      r2891 := rewire_littleendian_2736(r2890);
      null;
      null;
      null;
      null;
      r2893 := (r2619 & r2620 & r2621 & r2622);
      r2894 := rewire_littleendian_2736(r2893);
      null;
      null;
      null;
      null;
      r2896 := (r2623 & r2624 & r2625 & r2626);
      r2897 := rewire_littleendian_2736(r2896);
      null;
      null;
      null;
      null;
      r2899 := (r2627 & r2628 & r2629 & r2630);
      r2900 := rewire_littleendian_2736(r2899);
      null;
      null;
      null;
      null;
      r2902 := (r2631 & r2632 & r2633 & r2634);
      r2903 := rewire_littleendian_2736(r2902);
      null;
      null;
      null;
      null;
      r2905 := (r2635 & r2636 & r2637 & r2638);
      r2906 := rewire_littleendian_2736(r2905);
      null;
      null;
      null;
      null;
      r2908 := (r2639 & r2640 & r2641 & r2642);
      r2909 := rewire_littleendian_2736(r2908);
      null;
      null;
      null;
      null;
      r2911 := (r2643 & r2644 & r2645 & r2646);
      r2912 := rewire_littleendian_2736(r2911);
      null;
      null;
      null;
      null;
      r2914 := (r2647 & r2648 & r2649 & r2650);
      r2915 := rewire_littleendian_2736(r2914);
      null;
      null;
      null;
      null;
      r2917 := (r2651 & r2652 & r2653 & r2654);
      r2918 := rewire_littleendian_2736(r2917);
      null;
      null;
      null;
      null;
      r2920 := (r2655 & r2656 & r2657 & r2658);
      r2921 := rewire_littleendian_2736(r2920);
      null;
      null;
      null;
      null;
      r2923 := (r2659 & r2660 & r2661 & r2662);
      r2924 := rewire_littleendian_2736(r2923);
      null;
      null;
      null;
      null;
      r2926 := (r2663 & r2664 & r2665 & r2666);
      r2927 := rewire_littleendian_2736(r2926);
      null;
      null;
      null;
      null;
      r2929 := (r2667 & r2668 & r2669 & r2670);
      r2930 := rewire_littleendian_2736(r2929);
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      r2932 := (r2885 & r2888 & r2891 & r2894 & r2897 & r2900 & r2903 & r2906 & r2909 & r2912 & r2915 & r2918 & r2921 & r2924 & r2927 & r2930);
      r2605 := r2932;
    end if;
    return r2605;
  end rewire_impwords_2602;
  function rewire_littleendian_2736(r2737 : std_logic_vector) return std_logic_vector
  is
    variable r2882 : std_logic_vector(0 to 31) := (others => '0');
    variable r2881 : std_logic_vector(0 to 15) := (others => '0');
    variable r2880 : std_logic_vector(0 to 15) := (others => '0');
    variable r2834 : std_logic_vector(0 to 15) := (others => '0');
    variable r2833 : std_logic_vector(0 to 7) := (others => '0');
    variable r2832 : std_logic_vector(0 to 7) := (others => '0');
    variable r2753 : std_logic_vector(0 to 31) := (others => '0');
    variable r2752 : std_logic_vector(0 to 15) := (others => '0');
    variable r2751 : std_logic_vector(0 to 15) := (others => '0');
    variable b2749 : boolean := false;
    variable b2748 : boolean := false;
    variable b2747 : boolean := false;
    variable b2746 : boolean := false;
    variable b2745 : boolean := false;
    variable r2744 : std_logic_vector(0 to 7) := (others => '0');
    variable r2743 : std_logic_vector(0 to 7) := (others => '0');
    variable r2742 : std_logic_vector(0 to 7) := (others => '0');
    variable r2741 : std_logic_vector(0 to 7) := (others => '0');
    variable b2740 : boolean := false;
    variable r2739 : std_logic_vector(0 to 31) := (others => '0');
  begin
    b2740 := true;
    r2741 := r2737(0 to 7);
    r2742 := r2737(8 to 15);
    r2743 := r2737(16 to 23);
    r2744 := r2737(24 to 31);
    b2745 := true;
    b2746 := true;
    b2747 := true;
    b2748 := true;
    b2749 := (b2745 AND (b2746 AND (b2747 AND b2748)));
    if b2749 then
      null;
      null;
      r2880 := rewire_w8to16le_2831(r2744,r2743);
      null;
      null;
      r2881 := rewire_w8to16le_2831(r2742,r2741);
      r2882 := rewire_w16tow32le_2750(r2880,r2881);
      r2739 := r2882;
    end if;
    return r2739;
  end rewire_littleendian_2736;
  function rewire_w8to16le_2831(r2832 : std_logic_vector ; r2833 : std_logic_vector) return std_logic_vector
  is
    variable r2879 : std_logic_vector(0 to 15) := (others => '0');
    variable b2877 : boolean := false;
    variable b2876 : boolean := false;
    variable b2875 : boolean := false;
    variable b2874 : boolean := false;
    variable b2873 : boolean := false;
    variable b2872 : boolean := false;
    variable b2871 : boolean := false;
    variable b2870 : boolean := false;
    variable b2869 : boolean := false;
    variable b2868 : boolean := false;
    variable r2867 : std_logic_vector(0 to 0) := (others => '0');
    variable r2866 : std_logic_vector(0 to 0) := (others => '0');
    variable r2865 : std_logic_vector(0 to 0) := (others => '0');
    variable r2864 : std_logic_vector(0 to 0) := (others => '0');
    variable r2863 : std_logic_vector(0 to 0) := (others => '0');
    variable r2862 : std_logic_vector(0 to 0) := (others => '0');
    variable r2861 : std_logic_vector(0 to 0) := (others => '0');
    variable r2860 : std_logic_vector(0 to 0) := (others => '0');
    variable b2859 : boolean := false;
    variable b2858 : boolean := false;
    variable b2857 : boolean := false;
    variable b2856 : boolean := false;
    variable b2855 : boolean := false;
    variable b2854 : boolean := false;
    variable b2853 : boolean := false;
    variable b2852 : boolean := false;
    variable b2851 : boolean := false;
    variable b2850 : boolean := false;
    variable r2849 : std_logic_vector(0 to 0) := (others => '0');
    variable r2848 : std_logic_vector(0 to 0) := (others => '0');
    variable r2847 : std_logic_vector(0 to 0) := (others => '0');
    variable r2846 : std_logic_vector(0 to 0) := (others => '0');
    variable r2845 : std_logic_vector(0 to 0) := (others => '0');
    variable r2844 : std_logic_vector(0 to 0) := (others => '0');
    variable r2843 : std_logic_vector(0 to 0) := (others => '0');
    variable r2842 : std_logic_vector(0 to 0) := (others => '0');
    variable b2841 : boolean := false;
    variable r2840 : std_logic_vector(0 to 7) := (others => '0');
    variable r2839 : std_logic_vector(0 to 7) := (others => '0');
    variable b2838 : boolean := false;
    variable r2837 : std_logic_vector(0 to 15) := (others => '0');
    variable r2836 : std_logic_vector(0 to 15) := (others => '0');
  begin
    b2838 := true;
    r2839 := r2836(0 to 7);
    r2840 := r2836(8 to 15);
    b2841 := true;
    r2842 := r2839(0 to 0);
    r2843 := r2839(1 to 1);
    r2844 := r2839(2 to 2);
    r2845 := r2839(3 to 3);
    r2846 := r2839(4 to 4);
    r2847 := r2839(5 to 5);
    r2848 := r2839(6 to 6);
    r2849 := r2839(7 to 7);
    b2850 := true;
    b2851 := true;
    b2852 := true;
    b2853 := true;
    b2854 := true;
    b2855 := true;
    b2856 := true;
    b2857 := true;
    b2858 := (b2850 AND (b2851 AND (b2852 AND (b2853 AND (b2854 AND (b2855 AND (b2856 AND b2857)))))));
    b2859 := true;
    r2860 := r2840(0 to 0);
    r2861 := r2840(1 to 1);
    r2862 := r2840(2 to 2);
    r2863 := r2840(3 to 3);
    r2864 := r2840(4 to 4);
    r2865 := r2840(5 to 5);
    r2866 := r2840(6 to 6);
    r2867 := r2840(7 to 7);
    b2868 := true;
    b2869 := true;
    b2870 := true;
    b2871 := true;
    b2872 := true;
    b2873 := true;
    b2874 := true;
    b2875 := true;
    b2876 := (b2868 AND (b2869 AND (b2870 AND (b2871 AND (b2872 AND (b2873 AND (b2874 AND b2875)))))));
    b2877 := (b2858 AND b2876);
    if b2877 then
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      r2879 := (r2860 & r2861 & r2862 & r2863 & r2864 & r2865 & r2866 & r2867 & r2842 & r2843 & r2844 & r2845 & r2846 & r2847 & r2848 & r2849);
      r2837 := r2879;
    end if;
    return r2837;
  end rewire_w8to16le_2831;
  function rewire_w16tow32le_2750(r2751 : std_logic_vector ; r2752 : std_logic_vector) return std_logic_vector
  is
    variable r2830 : std_logic_vector(0 to 31) := (others => '0');
    variable b2828 : boolean := false;
    variable b2827 : boolean := false;
    variable b2826 : boolean := false;
    variable b2825 : boolean := false;
    variable b2824 : boolean := false;
    variable b2823 : boolean := false;
    variable b2822 : boolean := false;
    variable b2821 : boolean := false;
    variable b2820 : boolean := false;
    variable b2819 : boolean := false;
    variable b2818 : boolean := false;
    variable b2817 : boolean := false;
    variable b2816 : boolean := false;
    variable b2815 : boolean := false;
    variable b2814 : boolean := false;
    variable b2813 : boolean := false;
    variable b2812 : boolean := false;
    variable b2811 : boolean := false;
    variable r2810 : std_logic_vector(0 to 0) := (others => '0');
    variable r2809 : std_logic_vector(0 to 0) := (others => '0');
    variable r2808 : std_logic_vector(0 to 0) := (others => '0');
    variable r2807 : std_logic_vector(0 to 0) := (others => '0');
    variable r2806 : std_logic_vector(0 to 0) := (others => '0');
    variable r2805 : std_logic_vector(0 to 0) := (others => '0');
    variable r2804 : std_logic_vector(0 to 0) := (others => '0');
    variable r2803 : std_logic_vector(0 to 0) := (others => '0');
    variable r2802 : std_logic_vector(0 to 0) := (others => '0');
    variable r2801 : std_logic_vector(0 to 0) := (others => '0');
    variable r2800 : std_logic_vector(0 to 0) := (others => '0');
    variable r2799 : std_logic_vector(0 to 0) := (others => '0');
    variable r2798 : std_logic_vector(0 to 0) := (others => '0');
    variable r2797 : std_logic_vector(0 to 0) := (others => '0');
    variable r2796 : std_logic_vector(0 to 0) := (others => '0');
    variable r2795 : std_logic_vector(0 to 0) := (others => '0');
    variable b2794 : boolean := false;
    variable b2793 : boolean := false;
    variable b2792 : boolean := false;
    variable b2791 : boolean := false;
    variable b2790 : boolean := false;
    variable b2789 : boolean := false;
    variable b2788 : boolean := false;
    variable b2787 : boolean := false;
    variable b2786 : boolean := false;
    variable b2785 : boolean := false;
    variable b2784 : boolean := false;
    variable b2783 : boolean := false;
    variable b2782 : boolean := false;
    variable b2781 : boolean := false;
    variable b2780 : boolean := false;
    variable b2779 : boolean := false;
    variable b2778 : boolean := false;
    variable b2777 : boolean := false;
    variable r2776 : std_logic_vector(0 to 0) := (others => '0');
    variable r2775 : std_logic_vector(0 to 0) := (others => '0');
    variable r2774 : std_logic_vector(0 to 0) := (others => '0');
    variable r2773 : std_logic_vector(0 to 0) := (others => '0');
    variable r2772 : std_logic_vector(0 to 0) := (others => '0');
    variable r2771 : std_logic_vector(0 to 0) := (others => '0');
    variable r2770 : std_logic_vector(0 to 0) := (others => '0');
    variable r2769 : std_logic_vector(0 to 0) := (others => '0');
    variable r2768 : std_logic_vector(0 to 0) := (others => '0');
    variable r2767 : std_logic_vector(0 to 0) := (others => '0');
    variable r2766 : std_logic_vector(0 to 0) := (others => '0');
    variable r2765 : std_logic_vector(0 to 0) := (others => '0');
    variable r2764 : std_logic_vector(0 to 0) := (others => '0');
    variable r2763 : std_logic_vector(0 to 0) := (others => '0');
    variable r2762 : std_logic_vector(0 to 0) := (others => '0');
    variable r2761 : std_logic_vector(0 to 0) := (others => '0');
    variable b2760 : boolean := false;
    variable r2759 : std_logic_vector(0 to 15) := (others => '0');
    variable r2758 : std_logic_vector(0 to 15) := (others => '0');
    variable b2757 : boolean := false;
    variable r2756 : std_logic_vector(0 to 31) := (others => '0');
    variable r2755 : std_logic_vector(0 to 31) := (others => '0');
  begin
    b2757 := true;
    r2758 := r2755(0 to 15);
    r2759 := r2755(16 to 31);
    b2760 := true;
    r2761 := r2758(0 to 0);
    r2762 := r2758(1 to 1);
    r2763 := r2758(2 to 2);
    r2764 := r2758(3 to 3);
    r2765 := r2758(4 to 4);
    r2766 := r2758(5 to 5);
    r2767 := r2758(6 to 6);
    r2768 := r2758(7 to 7);
    r2769 := r2758(8 to 8);
    r2770 := r2758(9 to 9);
    r2771 := r2758(10 to 10);
    r2772 := r2758(11 to 11);
    r2773 := r2758(12 to 12);
    r2774 := r2758(13 to 13);
    r2775 := r2758(14 to 14);
    r2776 := r2758(15 to 15);
    b2777 := true;
    b2778 := true;
    b2779 := true;
    b2780 := true;
    b2781 := true;
    b2782 := true;
    b2783 := true;
    b2784 := true;
    b2785 := true;
    b2786 := true;
    b2787 := true;
    b2788 := true;
    b2789 := true;
    b2790 := true;
    b2791 := true;
    b2792 := true;
    b2793 := (b2777 AND (b2778 AND (b2779 AND (b2780 AND (b2781 AND (b2782 AND (b2783 AND (b2784 AND (b2785 AND (b2786 AND (b2787 AND (b2788 AND (b2789 AND (b2790 AND (b2791 AND b2792)))))))))))))));
    b2794 := true;
    r2795 := r2759(0 to 0);
    r2796 := r2759(1 to 1);
    r2797 := r2759(2 to 2);
    r2798 := r2759(3 to 3);
    r2799 := r2759(4 to 4);
    r2800 := r2759(5 to 5);
    r2801 := r2759(6 to 6);
    r2802 := r2759(7 to 7);
    r2803 := r2759(8 to 8);
    r2804 := r2759(9 to 9);
    r2805 := r2759(10 to 10);
    r2806 := r2759(11 to 11);
    r2807 := r2759(12 to 12);
    r2808 := r2759(13 to 13);
    r2809 := r2759(14 to 14);
    r2810 := r2759(15 to 15);
    b2811 := true;
    b2812 := true;
    b2813 := true;
    b2814 := true;
    b2815 := true;
    b2816 := true;
    b2817 := true;
    b2818 := true;
    b2819 := true;
    b2820 := true;
    b2821 := true;
    b2822 := true;
    b2823 := true;
    b2824 := true;
    b2825 := true;
    b2826 := true;
    b2827 := (b2811 AND (b2812 AND (b2813 AND (b2814 AND (b2815 AND (b2816 AND (b2817 AND (b2818 AND (b2819 AND (b2820 AND (b2821 AND (b2822 AND (b2823 AND (b2824 AND (b2825 AND b2826)))))))))))))));
    b2828 := (b2793 AND b2827);
    if b2828 then
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      r2830 := (r2761 & r2762 & r2763 & r2764 & r2765 & r2766 & r2767 & r2768 & r2769 & r2770 & r2771 & r2772 & r2773 & r2774 & r2775 & r2776 & r2795 & r2796 & r2797 & r2798 & r2799 & r2800 & r2801 & r2802 & r2803 & r2804 & r2805 & r2806 & r2807 & r2808 & r2809 & r2810);
      r2756 := r2830;
    end if;
    return r2756;
  end rewire_w16tow32le_2750;
  function rewire_salsaHashp_1978(r1979 : std_logic_vector) return std_logic_vector
  is
    variable r2601 : std_logic_vector(0 to 511) := (others => '0');
    variable r2600 : std_logic_vector(0 to 31) := (others => '0');
    variable r2599 : std_logic_vector(0 to 31) := (others => '0');
    variable r2598 : std_logic_vector(0 to 31) := (others => '0');
    variable r2597 : std_logic_vector(0 to 31) := (others => '0');
    variable r2596 : std_logic_vector(0 to 31) := (others => '0');
    variable r2595 : std_logic_vector(0 to 31) := (others => '0');
    variable r2594 : std_logic_vector(0 to 31) := (others => '0');
    variable r2593 : std_logic_vector(0 to 31) := (others => '0');
    variable r2592 : std_logic_vector(0 to 31) := (others => '0');
    variable r2591 : std_logic_vector(0 to 31) := (others => '0');
    variable r2590 : std_logic_vector(0 to 31) := (others => '0');
    variable r2589 : std_logic_vector(0 to 31) := (others => '0');
    variable r2588 : std_logic_vector(0 to 31) := (others => '0');
    variable r2587 : std_logic_vector(0 to 31) := (others => '0');
    variable r2586 : std_logic_vector(0 to 31) := (others => '0');
    variable r2585 : std_logic_vector(0 to 31) := (others => '0');
    variable b2583 : boolean := false;
    variable b2582 : boolean := false;
    variable b2581 : boolean := false;
    variable b2580 : boolean := false;
    variable b2579 : boolean := false;
    variable b2578 : boolean := false;
    variable b2577 : boolean := false;
    variable b2576 : boolean := false;
    variable b2575 : boolean := false;
    variable b2574 : boolean := false;
    variable b2573 : boolean := false;
    variable b2572 : boolean := false;
    variable b2571 : boolean := false;
    variable b2570 : boolean := false;
    variable b2569 : boolean := false;
    variable b2568 : boolean := false;
    variable b2567 : boolean := false;
    variable r2566 : std_logic_vector(0 to 31) := (others => '0');
    variable r2565 : std_logic_vector(0 to 31) := (others => '0');
    variable r2564 : std_logic_vector(0 to 31) := (others => '0');
    variable r2563 : std_logic_vector(0 to 31) := (others => '0');
    variable r2562 : std_logic_vector(0 to 31) := (others => '0');
    variable r2561 : std_logic_vector(0 to 31) := (others => '0');
    variable r2560 : std_logic_vector(0 to 31) := (others => '0');
    variable r2559 : std_logic_vector(0 to 31) := (others => '0');
    variable r2558 : std_logic_vector(0 to 31) := (others => '0');
    variable r2557 : std_logic_vector(0 to 31) := (others => '0');
    variable r2556 : std_logic_vector(0 to 31) := (others => '0');
    variable r2555 : std_logic_vector(0 to 31) := (others => '0');
    variable r2554 : std_logic_vector(0 to 31) := (others => '0');
    variable r2553 : std_logic_vector(0 to 31) := (others => '0');
    variable r2552 : std_logic_vector(0 to 31) := (others => '0');
    variable r2551 : std_logic_vector(0 to 31) := (others => '0');
    variable b2550 : boolean := false;
    variable r2549 : std_logic_vector(0 to 511) := (others => '0');
    variable r2548 : std_logic_vector(0 to 511) := (others => '0');
    variable r2547 : std_logic_vector(0 to 511) := (others => '0');
    variable r2546 : std_logic_vector(0 to 511) := (others => '0');
    variable r2545 : std_logic_vector(0 to 511) := (others => '0');
    variable r2544 : std_logic_vector(0 to 511) := (others => '0');
    variable r2543 : std_logic_vector(0 to 511) := (others => '0');
    variable r2542 : std_logic_vector(0 to 511) := (others => '0');
    variable r2541 : std_logic_vector(0 to 511) := (others => '0');
    variable r2540 : std_logic_vector(0 to 511) := (others => '0');
    variable r2539 : std_logic_vector(0 to 511) := (others => '0');
    variable r2018 : std_logic_vector(0 to 511) := (others => '0');
    variable r2017 : std_logic_vector(0 to 511) := (others => '0');
    variable b2015 : boolean := false;
    variable b2014 : boolean := false;
    variable b2013 : boolean := false;
    variable b2012 : boolean := false;
    variable b2011 : boolean := false;
    variable b2010 : boolean := false;
    variable b2009 : boolean := false;
    variable b2008 : boolean := false;
    variable b2007 : boolean := false;
    variable b2006 : boolean := false;
    variable b2005 : boolean := false;
    variable b2004 : boolean := false;
    variable b2003 : boolean := false;
    variable b2002 : boolean := false;
    variable b2001 : boolean := false;
    variable b2000 : boolean := false;
    variable b1999 : boolean := false;
    variable r1998 : std_logic_vector(0 to 31) := (others => '0');
    variable r1997 : std_logic_vector(0 to 31) := (others => '0');
    variable r1996 : std_logic_vector(0 to 31) := (others => '0');
    variable r1995 : std_logic_vector(0 to 31) := (others => '0');
    variable r1994 : std_logic_vector(0 to 31) := (others => '0');
    variable r1993 : std_logic_vector(0 to 31) := (others => '0');
    variable r1992 : std_logic_vector(0 to 31) := (others => '0');
    variable r1991 : std_logic_vector(0 to 31) := (others => '0');
    variable r1990 : std_logic_vector(0 to 31) := (others => '0');
    variable r1989 : std_logic_vector(0 to 31) := (others => '0');
    variable r1988 : std_logic_vector(0 to 31) := (others => '0');
    variable r1987 : std_logic_vector(0 to 31) := (others => '0');
    variable r1986 : std_logic_vector(0 to 31) := (others => '0');
    variable r1985 : std_logic_vector(0 to 31) := (others => '0');
    variable r1984 : std_logic_vector(0 to 31) := (others => '0');
    variable r1983 : std_logic_vector(0 to 31) := (others => '0');
    variable b1982 : boolean := false;
    variable r1981 : std_logic_vector(0 to 511) := (others => '0');
  begin
    b1982 := true;
    r1983 := r1979(0 to 31);
    r1984 := r1979(32 to 63);
    r1985 := r1979(64 to 95);
    r1986 := r1979(96 to 127);
    r1987 := r1979(128 to 159);
    r1988 := r1979(160 to 191);
    r1989 := r1979(192 to 223);
    r1990 := r1979(224 to 255);
    r1991 := r1979(256 to 287);
    r1992 := r1979(288 to 319);
    r1993 := r1979(320 to 351);
    r1994 := r1979(352 to 383);
    r1995 := r1979(384 to 415);
    r1996 := r1979(416 to 447);
    r1997 := r1979(448 to 479);
    r1998 := r1979(480 to 511);
    b1999 := true;
    b2000 := true;
    b2001 := true;
    b2002 := true;
    b2003 := true;
    b2004 := true;
    b2005 := true;
    b2006 := true;
    b2007 := true;
    b2008 := true;
    b2009 := true;
    b2010 := true;
    b2011 := true;
    b2012 := true;
    b2013 := true;
    b2014 := true;
    b2015 := (b1999 AND (b2000 AND (b2001 AND (b2002 AND (b2003 AND (b2004 AND (b2005 AND (b2006 AND (b2007 AND (b2008 AND (b2009 AND (b2010 AND (b2011 AND (b2012 AND (b2013 AND b2014)))))))))))))));
    if b2015 then
      b2550 := true;
      r2551 := r2548(0 to 31);
      r2552 := r2548(32 to 63);
      r2553 := r2548(64 to 95);
      r2554 := r2548(96 to 127);
      r2555 := r2548(128 to 159);
      r2556 := r2548(160 to 191);
      r2557 := r2548(192 to 223);
      r2558 := r2548(224 to 255);
      r2559 := r2548(256 to 287);
      r2560 := r2548(288 to 319);
      r2561 := r2548(320 to 351);
      r2562 := r2548(352 to 383);
      r2563 := r2548(384 to 415);
      r2564 := r2548(416 to 447);
      r2565 := r2548(448 to 479);
      r2566 := r2548(480 to 511);
      b2567 := true;
      b2568 := true;
      b2569 := true;
      b2570 := true;
      b2571 := true;
      b2572 := true;
      b2573 := true;
      b2574 := true;
      b2575 := true;
      b2576 := true;
      b2577 := true;
      b2578 := true;
      b2579 := true;
      b2580 := true;
      b2581 := true;
      b2582 := true;
      b2583 := (b2567 AND (b2568 AND (b2569 AND (b2570 AND (b2571 AND (b2572 AND (b2573 AND (b2574 AND (b2575 AND (b2576 AND (b2577 AND (b2578 AND (b2579 AND (b2580 AND (b2581 AND b2582)))))))))))))));
      if b2583 then
        null;
        null;
        r2585 := add32(r2551,r1983);
        null;
        null;
        r2586 := add32(r2552,r1984);
        null;
        null;
        r2587 := add32(r2553,r1985);
        null;
        null;
        r2588 := add32(r2554,r1986);
        null;
        null;
        r2589 := add32(r2555,r1987);
        null;
        null;
        r2590 := add32(r2556,r1988);
        null;
        null;
        r2591 := add32(r2557,r1989);
        null;
        null;
        r2592 := add32(r2558,r1990);
        null;
        null;
        r2593 := add32(r2559,r1991);
        null;
        null;
        r2594 := add32(r2560,r1992);
        null;
        null;
        r2595 := add32(r2561,r1993);
        null;
        null;
        r2596 := add32(r2562,r1994);
        null;
        null;
        r2597 := add32(r2563,r1995);
        null;
        null;
        r2598 := add32(r2564,r1996);
        null;
        null;
        r2599 := add32(r2565,r1997);
        null;
        null;
        r2600 := add32(r2566,r1998);
        r2601 := (r2585 & r2586 & r2587 & r2588 & r2589 & r2590 & r2591 & r2592 & r2593 & r2594 & r2595 & r2596 & r2597 & r2598 & r2599 & r2600);
        r2549 := r2601;
      end if;
      r1981 := r2549;
    end if;
    return r1981;
  end rewire_salsaHashp_1978;
  function rewire_doubleRound_2016(r2017 : std_logic_vector) return std_logic_vector
  is
    variable r2538 : std_logic_vector(0 to 511) := (others => '0');
    variable r2537 : std_logic_vector(0 to 511) := (others => '0');
    variable r2438 : std_logic_vector(0 to 511) := (others => '0');
    variable r2437 : std_logic_vector(0 to 511) := (others => '0');
    variable r2021 : std_logic_vector(0 to 511) := (others => '0');
    variable r2020 : std_logic_vector(0 to 511) := (others => '0');
  begin
    null;
    r2537 := rewire_columnRound_2436(r2017);
    r2538 := rewire_rowRound_2019(r2537);
    return r2538;
  end rewire_doubleRound_2016;
  function rewire_columnRound_2436(r2437 : std_logic_vector) return std_logic_vector
  is
    variable r2536 : std_logic_vector(0 to 511) := (others => '0');
    variable b2534 : boolean := false;
    variable b2533 : boolean := false;
    variable b2532 : boolean := false;
    variable b2531 : boolean := false;
    variable b2530 : boolean := false;
    variable b2529 : boolean := false;
    variable r2528 : std_logic_vector(0 to 31) := (others => '0');
    variable r2527 : std_logic_vector(0 to 31) := (others => '0');
    variable r2526 : std_logic_vector(0 to 31) := (others => '0');
    variable r2525 : std_logic_vector(0 to 31) := (others => '0');
    variable b2524 : boolean := false;
    variable b2523 : boolean := false;
    variable b2522 : boolean := false;
    variable b2521 : boolean := false;
    variable b2520 : boolean := false;
    variable b2519 : boolean := false;
    variable r2518 : std_logic_vector(0 to 31) := (others => '0');
    variable r2517 : std_logic_vector(0 to 31) := (others => '0');
    variable r2516 : std_logic_vector(0 to 31) := (others => '0');
    variable r2515 : std_logic_vector(0 to 31) := (others => '0');
    variable b2514 : boolean := false;
    variable b2513 : boolean := false;
    variable b2512 : boolean := false;
    variable b2511 : boolean := false;
    variable b2510 : boolean := false;
    variable b2509 : boolean := false;
    variable r2508 : std_logic_vector(0 to 31) := (others => '0');
    variable r2507 : std_logic_vector(0 to 31) := (others => '0');
    variable r2506 : std_logic_vector(0 to 31) := (others => '0');
    variable r2505 : std_logic_vector(0 to 31) := (others => '0');
    variable b2504 : boolean := false;
    variable b2503 : boolean := false;
    variable b2502 : boolean := false;
    variable b2501 : boolean := false;
    variable b2500 : boolean := false;
    variable b2499 : boolean := false;
    variable r2498 : std_logic_vector(0 to 31) := (others => '0');
    variable r2497 : std_logic_vector(0 to 31) := (others => '0');
    variable r2496 : std_logic_vector(0 to 31) := (others => '0');
    variable r2495 : std_logic_vector(0 to 31) := (others => '0');
    variable b2494 : boolean := false;
    variable r2493 : std_logic_vector(0 to 127) := (others => '0');
    variable r2492 : std_logic_vector(0 to 127) := (others => '0');
    variable r2491 : std_logic_vector(0 to 127) := (others => '0');
    variable r2490 : std_logic_vector(0 to 127) := (others => '0');
    variable b2489 : boolean := false;
    variable r2488 : std_logic_vector(0 to 511) := (others => '0');
    variable r2487 : std_logic_vector(0 to 511) := (others => '0');
    variable r2485 : std_logic_vector(0 to 127) := (others => '0');
    variable r2484 : std_logic_vector(0 to 127) := (others => '0');
    variable r2482 : std_logic_vector(0 to 127) := (others => '0');
    variable r2481 : std_logic_vector(0 to 127) := (others => '0');
    variable r2479 : std_logic_vector(0 to 127) := (others => '0');
    variable r2478 : std_logic_vector(0 to 127) := (others => '0');
    variable r2476 : std_logic_vector(0 to 127) := (others => '0');
    variable r2475 : std_logic_vector(0 to 127) := (others => '0');
    variable b2473 : boolean := false;
    variable b2472 : boolean := false;
    variable b2471 : boolean := false;
    variable b2470 : boolean := false;
    variable b2469 : boolean := false;
    variable b2468 : boolean := false;
    variable b2467 : boolean := false;
    variable b2466 : boolean := false;
    variable b2465 : boolean := false;
    variable b2464 : boolean := false;
    variable b2463 : boolean := false;
    variable b2462 : boolean := false;
    variable b2461 : boolean := false;
    variable b2460 : boolean := false;
    variable b2459 : boolean := false;
    variable b2458 : boolean := false;
    variable b2457 : boolean := false;
    variable r2456 : std_logic_vector(0 to 31) := (others => '0');
    variable r2455 : std_logic_vector(0 to 31) := (others => '0');
    variable r2454 : std_logic_vector(0 to 31) := (others => '0');
    variable r2453 : std_logic_vector(0 to 31) := (others => '0');
    variable r2452 : std_logic_vector(0 to 31) := (others => '0');
    variable r2451 : std_logic_vector(0 to 31) := (others => '0');
    variable r2450 : std_logic_vector(0 to 31) := (others => '0');
    variable r2449 : std_logic_vector(0 to 31) := (others => '0');
    variable r2448 : std_logic_vector(0 to 31) := (others => '0');
    variable r2447 : std_logic_vector(0 to 31) := (others => '0');
    variable r2446 : std_logic_vector(0 to 31) := (others => '0');
    variable r2445 : std_logic_vector(0 to 31) := (others => '0');
    variable r2444 : std_logic_vector(0 to 31) := (others => '0');
    variable r2443 : std_logic_vector(0 to 31) := (others => '0');
    variable r2442 : std_logic_vector(0 to 31) := (others => '0');
    variable r2441 : std_logic_vector(0 to 31) := (others => '0');
    variable b2440 : boolean := false;
    variable r2439 : std_logic_vector(0 to 511) := (others => '0');
  begin
    b2440 := true;
    r2441 := r2437(0 to 31);
    r2442 := r2437(32 to 63);
    r2443 := r2437(64 to 95);
    r2444 := r2437(96 to 127);
    r2445 := r2437(128 to 159);
    r2446 := r2437(160 to 191);
    r2447 := r2437(192 to 223);
    r2448 := r2437(224 to 255);
    r2449 := r2437(256 to 287);
    r2450 := r2437(288 to 319);
    r2451 := r2437(320 to 351);
    r2452 := r2437(352 to 383);
    r2453 := r2437(384 to 415);
    r2454 := r2437(416 to 447);
    r2455 := r2437(448 to 479);
    r2456 := r2437(480 to 511);
    b2457 := true;
    b2458 := true;
    b2459 := true;
    b2460 := true;
    b2461 := true;
    b2462 := true;
    b2463 := true;
    b2464 := true;
    b2465 := true;
    b2466 := true;
    b2467 := true;
    b2468 := true;
    b2469 := true;
    b2470 := true;
    b2471 := true;
    b2472 := true;
    b2473 := (b2457 AND (b2458 AND (b2459 AND (b2460 AND (b2461 AND (b2462 AND (b2463 AND (b2464 AND (b2465 AND (b2466 AND (b2467 AND (b2468 AND (b2469 AND (b2470 AND (b2471 AND b2472)))))))))))))));
    if b2473 then
      null;
      null;
      null;
      null;
      r2475 := (r2441 & r2445 & r2449 & r2453);
      r2476 := rewire_quarterRound_2057(r2475);
      null;
      null;
      null;
      null;
      r2478 := (r2446 & r2450 & r2454 & r2442);
      r2479 := rewire_quarterRound_2057(r2478);
      null;
      null;
      null;
      null;
      r2481 := (r2451 & r2455 & r2443 & r2447);
      r2482 := rewire_quarterRound_2057(r2481);
      null;
      null;
      null;
      null;
      r2484 := (r2456 & r2444 & r2448 & r2452);
      r2485 := rewire_quarterRound_2057(r2484);
      b2489 := true;
      r2490 := r2487(0 to 127);
      r2491 := r2487(128 to 255);
      r2492 := r2487(256 to 383);
      r2493 := r2487(384 to 511);
      b2494 := true;
      r2495 := r2490(0 to 31);
      r2496 := r2490(32 to 63);
      r2497 := r2490(64 to 95);
      r2498 := r2490(96 to 127);
      b2499 := true;
      b2500 := true;
      b2501 := true;
      b2502 := true;
      b2503 := (b2499 AND (b2500 AND (b2501 AND b2502)));
      b2504 := true;
      r2505 := r2491(0 to 31);
      r2506 := r2491(32 to 63);
      r2507 := r2491(64 to 95);
      r2508 := r2491(96 to 127);
      b2509 := true;
      b2510 := true;
      b2511 := true;
      b2512 := true;
      b2513 := (b2509 AND (b2510 AND (b2511 AND b2512)));
      b2514 := true;
      r2515 := r2492(0 to 31);
      r2516 := r2492(32 to 63);
      r2517 := r2492(64 to 95);
      r2518 := r2492(96 to 127);
      b2519 := true;
      b2520 := true;
      b2521 := true;
      b2522 := true;
      b2523 := (b2519 AND (b2520 AND (b2521 AND b2522)));
      b2524 := true;
      r2525 := r2493(0 to 31);
      r2526 := r2493(32 to 63);
      r2527 := r2493(64 to 95);
      r2528 := r2493(96 to 127);
      b2529 := true;
      b2530 := true;
      b2531 := true;
      b2532 := true;
      b2533 := (b2529 AND (b2530 AND (b2531 AND b2532)));
      b2534 := (b2503 AND (b2513 AND (b2523 AND b2533)));
      if b2534 then
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        r2536 := (r2495 & r2508 & r2517 & r2526 & r2496 & r2505 & r2518 & r2527 & r2497 & r2506 & r2515 & r2528 & r2498 & r2507 & r2516 & r2525);
        r2488 := r2536;
      end if;
      r2439 := r2488;
    end if;
    return r2439;
  end rewire_columnRound_2436;
  function rewire_rowRound_2019(r2020 : std_logic_vector) return std_logic_vector
  is
    variable r2435 : std_logic_vector(0 to 511) := (others => '0');
    variable b2433 : boolean := false;
    variable b2432 : boolean := false;
    variable b2431 : boolean := false;
    variable b2430 : boolean := false;
    variable b2429 : boolean := false;
    variable b2428 : boolean := false;
    variable r2427 : std_logic_vector(0 to 31) := (others => '0');
    variable r2426 : std_logic_vector(0 to 31) := (others => '0');
    variable r2425 : std_logic_vector(0 to 31) := (others => '0');
    variable r2424 : std_logic_vector(0 to 31) := (others => '0');
    variable b2423 : boolean := false;
    variable b2422 : boolean := false;
    variable b2421 : boolean := false;
    variable b2420 : boolean := false;
    variable b2419 : boolean := false;
    variable b2418 : boolean := false;
    variable r2417 : std_logic_vector(0 to 31) := (others => '0');
    variable r2416 : std_logic_vector(0 to 31) := (others => '0');
    variable r2415 : std_logic_vector(0 to 31) := (others => '0');
    variable r2414 : std_logic_vector(0 to 31) := (others => '0');
    variable b2413 : boolean := false;
    variable b2412 : boolean := false;
    variable b2411 : boolean := false;
    variable b2410 : boolean := false;
    variable b2409 : boolean := false;
    variable b2408 : boolean := false;
    variable r2407 : std_logic_vector(0 to 31) := (others => '0');
    variable r2406 : std_logic_vector(0 to 31) := (others => '0');
    variable r2405 : std_logic_vector(0 to 31) := (others => '0');
    variable r2404 : std_logic_vector(0 to 31) := (others => '0');
    variable b2403 : boolean := false;
    variable b2402 : boolean := false;
    variable b2401 : boolean := false;
    variable b2400 : boolean := false;
    variable b2399 : boolean := false;
    variable b2398 : boolean := false;
    variable r2397 : std_logic_vector(0 to 31) := (others => '0');
    variable r2396 : std_logic_vector(0 to 31) := (others => '0');
    variable r2395 : std_logic_vector(0 to 31) := (others => '0');
    variable r2394 : std_logic_vector(0 to 31) := (others => '0');
    variable b2393 : boolean := false;
    variable r2392 : std_logic_vector(0 to 127) := (others => '0');
    variable r2391 : std_logic_vector(0 to 127) := (others => '0');
    variable r2390 : std_logic_vector(0 to 127) := (others => '0');
    variable r2389 : std_logic_vector(0 to 127) := (others => '0');
    variable b2388 : boolean := false;
    variable r2387 : std_logic_vector(0 to 511) := (others => '0');
    variable r2386 : std_logic_vector(0 to 511) := (others => '0');
    variable r2384 : std_logic_vector(0 to 127) := (others => '0');
    variable r2383 : std_logic_vector(0 to 127) := (others => '0');
    variable r2381 : std_logic_vector(0 to 127) := (others => '0');
    variable r2380 : std_logic_vector(0 to 127) := (others => '0');
    variable r2378 : std_logic_vector(0 to 127) := (others => '0');
    variable r2377 : std_logic_vector(0 to 127) := (others => '0');
    variable r2375 : std_logic_vector(0 to 127) := (others => '0');
    variable r2374 : std_logic_vector(0 to 127) := (others => '0');
    variable r2059 : std_logic_vector(0 to 127) := (others => '0');
    variable r2058 : std_logic_vector(0 to 127) := (others => '0');
    variable b2056 : boolean := false;
    variable b2055 : boolean := false;
    variable b2054 : boolean := false;
    variable b2053 : boolean := false;
    variable b2052 : boolean := false;
    variable b2051 : boolean := false;
    variable b2050 : boolean := false;
    variable b2049 : boolean := false;
    variable b2048 : boolean := false;
    variable b2047 : boolean := false;
    variable b2046 : boolean := false;
    variable b2045 : boolean := false;
    variable b2044 : boolean := false;
    variable b2043 : boolean := false;
    variable b2042 : boolean := false;
    variable b2041 : boolean := false;
    variable b2040 : boolean := false;
    variable r2039 : std_logic_vector(0 to 31) := (others => '0');
    variable r2038 : std_logic_vector(0 to 31) := (others => '0');
    variable r2037 : std_logic_vector(0 to 31) := (others => '0');
    variable r2036 : std_logic_vector(0 to 31) := (others => '0');
    variable r2035 : std_logic_vector(0 to 31) := (others => '0');
    variable r2034 : std_logic_vector(0 to 31) := (others => '0');
    variable r2033 : std_logic_vector(0 to 31) := (others => '0');
    variable r2032 : std_logic_vector(0 to 31) := (others => '0');
    variable r2031 : std_logic_vector(0 to 31) := (others => '0');
    variable r2030 : std_logic_vector(0 to 31) := (others => '0');
    variable r2029 : std_logic_vector(0 to 31) := (others => '0');
    variable r2028 : std_logic_vector(0 to 31) := (others => '0');
    variable r2027 : std_logic_vector(0 to 31) := (others => '0');
    variable r2026 : std_logic_vector(0 to 31) := (others => '0');
    variable r2025 : std_logic_vector(0 to 31) := (others => '0');
    variable r2024 : std_logic_vector(0 to 31) := (others => '0');
    variable b2023 : boolean := false;
    variable r2022 : std_logic_vector(0 to 511) := (others => '0');
  begin
    b2023 := true;
    r2024 := r2020(0 to 31);
    r2025 := r2020(32 to 63);
    r2026 := r2020(64 to 95);
    r2027 := r2020(96 to 127);
    r2028 := r2020(128 to 159);
    r2029 := r2020(160 to 191);
    r2030 := r2020(192 to 223);
    r2031 := r2020(224 to 255);
    r2032 := r2020(256 to 287);
    r2033 := r2020(288 to 319);
    r2034 := r2020(320 to 351);
    r2035 := r2020(352 to 383);
    r2036 := r2020(384 to 415);
    r2037 := r2020(416 to 447);
    r2038 := r2020(448 to 479);
    r2039 := r2020(480 to 511);
    b2040 := true;
    b2041 := true;
    b2042 := true;
    b2043 := true;
    b2044 := true;
    b2045 := true;
    b2046 := true;
    b2047 := true;
    b2048 := true;
    b2049 := true;
    b2050 := true;
    b2051 := true;
    b2052 := true;
    b2053 := true;
    b2054 := true;
    b2055 := true;
    b2056 := (b2040 AND (b2041 AND (b2042 AND (b2043 AND (b2044 AND (b2045 AND (b2046 AND (b2047 AND (b2048 AND (b2049 AND (b2050 AND (b2051 AND (b2052 AND (b2053 AND (b2054 AND b2055)))))))))))))));
    if b2056 then
      null;
      null;
      null;
      null;
      r2374 := (r2024 & r2025 & r2026 & r2027);
      r2375 := rewire_quarterRound_2057(r2374);
      null;
      null;
      null;
      null;
      r2377 := (r2029 & r2030 & r2031 & r2028);
      r2378 := rewire_quarterRound_2057(r2377);
      null;
      null;
      null;
      null;
      r2380 := (r2034 & r2035 & r2032 & r2033);
      r2381 := rewire_quarterRound_2057(r2380);
      null;
      null;
      null;
      null;
      r2383 := (r2039 & r2036 & r2037 & r2038);
      r2384 := rewire_quarterRound_2057(r2383);
      b2388 := true;
      r2389 := r2386(0 to 127);
      r2390 := r2386(128 to 255);
      r2391 := r2386(256 to 383);
      r2392 := r2386(384 to 511);
      b2393 := true;
      r2394 := r2389(0 to 31);
      r2395 := r2389(32 to 63);
      r2396 := r2389(64 to 95);
      r2397 := r2389(96 to 127);
      b2398 := true;
      b2399 := true;
      b2400 := true;
      b2401 := true;
      b2402 := (b2398 AND (b2399 AND (b2400 AND b2401)));
      b2403 := true;
      r2404 := r2390(0 to 31);
      r2405 := r2390(32 to 63);
      r2406 := r2390(64 to 95);
      r2407 := r2390(96 to 127);
      b2408 := true;
      b2409 := true;
      b2410 := true;
      b2411 := true;
      b2412 := (b2408 AND (b2409 AND (b2410 AND b2411)));
      b2413 := true;
      r2414 := r2391(0 to 31);
      r2415 := r2391(32 to 63);
      r2416 := r2391(64 to 95);
      r2417 := r2391(96 to 127);
      b2418 := true;
      b2419 := true;
      b2420 := true;
      b2421 := true;
      b2422 := (b2418 AND (b2419 AND (b2420 AND b2421)));
      b2423 := true;
      r2424 := r2392(0 to 31);
      r2425 := r2392(32 to 63);
      r2426 := r2392(64 to 95);
      r2427 := r2392(96 to 127);
      b2428 := true;
      b2429 := true;
      b2430 := true;
      b2431 := true;
      b2432 := (b2428 AND (b2429 AND (b2430 AND b2431)));
      b2433 := (b2402 AND (b2412 AND (b2422 AND b2432)));
      if b2433 then
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        r2435 := (r2394 & r2395 & r2396 & r2397 & r2407 & r2404 & r2405 & r2406 & r2416 & r2417 & r2414 & r2415 & r2425 & r2426 & r2427 & r2424);
        r2387 := r2435;
      end if;
      r2022 := r2387;
    end if;
    return r2022;
  end rewire_rowRound_2019;
  function rewire_quarterRound_2057(r2058 : std_logic_vector) return std_logic_vector
  is
    variable r2372 : std_logic_vector(0 to 127) := (others => '0');
    variable r2370 : std_logic_vector(0 to 31) := (others => '0');
    variable r2369 : std_logic_vector(0 to 31) := (others => '0');
    variable r2368 : std_logic_vector(0 to 31) := (others => '0');
    variable r2298 : std_logic_vector(0 to 31) := (others => '0');
    variable r2297 : std_logic_vector(0 to 31) := (others => '0');
    variable r2295 : std_logic_vector(0 to 31) := (others => '0');
    variable r2294 : std_logic_vector(0 to 31) := (others => '0');
    variable r2293 : std_logic_vector(0 to 31) := (others => '0');
    variable r2223 : std_logic_vector(0 to 31) := (others => '0');
    variable r2222 : std_logic_vector(0 to 31) := (others => '0');
    variable r2220 : std_logic_vector(0 to 31) := (others => '0');
    variable r2219 : std_logic_vector(0 to 31) := (others => '0');
    variable r2218 : std_logic_vector(0 to 31) := (others => '0');
    variable r2148 : std_logic_vector(0 to 31) := (others => '0');
    variable r2147 : std_logic_vector(0 to 31) := (others => '0');
    variable r2145 : std_logic_vector(0 to 31) := (others => '0');
    variable r2144 : std_logic_vector(0 to 31) := (others => '0');
    variable r2143 : std_logic_vector(0 to 31) := (others => '0');
    variable r2073 : std_logic_vector(0 to 31) := (others => '0');
    variable r2072 : std_logic_vector(0 to 31) := (others => '0');
    variable b2070 : boolean := false;
    variable b2069 : boolean := false;
    variable b2068 : boolean := false;
    variable b2067 : boolean := false;
    variable b2066 : boolean := false;
    variable r2065 : std_logic_vector(0 to 31) := (others => '0');
    variable r2064 : std_logic_vector(0 to 31) := (others => '0');
    variable r2063 : std_logic_vector(0 to 31) := (others => '0');
    variable r2062 : std_logic_vector(0 to 31) := (others => '0');
    variable b2061 : boolean := false;
    variable r2060 : std_logic_vector(0 to 127) := (others => '0');
  begin
    b2061 := true;
    r2062 := r2058(0 to 31);
    r2063 := r2058(32 to 63);
    r2064 := r2058(64 to 95);
    r2065 := r2058(96 to 127);
    b2066 := true;
    b2067 := true;
    b2068 := true;
    b2069 := true;
    b2070 := (b2066 AND (b2067 AND (b2068 AND b2069)));
    if b2070 then
      null;
      null;
      null;
      r2143 := add32(r2062,r2065);
      r2144 := rewire_rot7_2071(r2143);
      r2145 := xor32(r2063,r2144);
      null;
      null;
      null;
      r2218 := add32(r2145,r2062);
      r2219 := rewire_rot9_2146(r2218);
      r2220 := xor32(r2064,r2219);
      null;
      null;
      null;
      r2293 := add32(r2220,r2145);
      r2294 := rewire_rot13_2221(r2293);
      r2295 := xor32(r2065,r2294);
      null;
      null;
      null;
      r2368 := add32(r2295,r2220);
      r2369 := rewire_rot18_2296(r2368);
      r2370 := xor32(r2062,r2369);
      null;
      null;
      null;
      null;
      r2372 := (r2370 & r2145 & r2220 & r2295);
      r2060 := r2372;
    end if;
    return r2060;
  end rewire_quarterRound_2057;
  function rewire_rot18_2296(r2297 : std_logic_vector) return std_logic_vector
  is
    variable r2367 : std_logic_vector(0 to 31) := (others => '0');
    variable b2365 : boolean := false;
    variable b2364 : boolean := false;
    variable b2363 : boolean := false;
    variable b2362 : boolean := false;
    variable b2361 : boolean := false;
    variable b2360 : boolean := false;
    variable b2359 : boolean := false;
    variable b2358 : boolean := false;
    variable b2357 : boolean := false;
    variable b2356 : boolean := false;
    variable b2355 : boolean := false;
    variable b2354 : boolean := false;
    variable b2353 : boolean := false;
    variable b2352 : boolean := false;
    variable b2351 : boolean := false;
    variable b2350 : boolean := false;
    variable b2349 : boolean := false;
    variable b2348 : boolean := false;
    variable b2347 : boolean := false;
    variable b2346 : boolean := false;
    variable b2345 : boolean := false;
    variable b2344 : boolean := false;
    variable b2343 : boolean := false;
    variable b2342 : boolean := false;
    variable b2341 : boolean := false;
    variable b2340 : boolean := false;
    variable b2339 : boolean := false;
    variable b2338 : boolean := false;
    variable b2337 : boolean := false;
    variable b2336 : boolean := false;
    variable b2335 : boolean := false;
    variable b2334 : boolean := false;
    variable b2333 : boolean := false;
    variable r2332 : std_logic_vector(0 to 0) := (others => '0');
    variable r2331 : std_logic_vector(0 to 0) := (others => '0');
    variable r2330 : std_logic_vector(0 to 0) := (others => '0');
    variable r2329 : std_logic_vector(0 to 0) := (others => '0');
    variable r2328 : std_logic_vector(0 to 0) := (others => '0');
    variable r2327 : std_logic_vector(0 to 0) := (others => '0');
    variable r2326 : std_logic_vector(0 to 0) := (others => '0');
    variable r2325 : std_logic_vector(0 to 0) := (others => '0');
    variable r2324 : std_logic_vector(0 to 0) := (others => '0');
    variable r2323 : std_logic_vector(0 to 0) := (others => '0');
    variable r2322 : std_logic_vector(0 to 0) := (others => '0');
    variable r2321 : std_logic_vector(0 to 0) := (others => '0');
    variable r2320 : std_logic_vector(0 to 0) := (others => '0');
    variable r2319 : std_logic_vector(0 to 0) := (others => '0');
    variable r2318 : std_logic_vector(0 to 0) := (others => '0');
    variable r2317 : std_logic_vector(0 to 0) := (others => '0');
    variable r2316 : std_logic_vector(0 to 0) := (others => '0');
    variable r2315 : std_logic_vector(0 to 0) := (others => '0');
    variable r2314 : std_logic_vector(0 to 0) := (others => '0');
    variable r2313 : std_logic_vector(0 to 0) := (others => '0');
    variable r2312 : std_logic_vector(0 to 0) := (others => '0');
    variable r2311 : std_logic_vector(0 to 0) := (others => '0');
    variable r2310 : std_logic_vector(0 to 0) := (others => '0');
    variable r2309 : std_logic_vector(0 to 0) := (others => '0');
    variable r2308 : std_logic_vector(0 to 0) := (others => '0');
    variable r2307 : std_logic_vector(0 to 0) := (others => '0');
    variable r2306 : std_logic_vector(0 to 0) := (others => '0');
    variable r2305 : std_logic_vector(0 to 0) := (others => '0');
    variable r2304 : std_logic_vector(0 to 0) := (others => '0');
    variable r2303 : std_logic_vector(0 to 0) := (others => '0');
    variable r2302 : std_logic_vector(0 to 0) := (others => '0');
    variable r2301 : std_logic_vector(0 to 0) := (others => '0');
    variable b2300 : boolean := false;
    variable r2299 : std_logic_vector(0 to 31) := (others => '0');
  begin
    b2300 := true;
    r2301 := r2297(0 to 0);
    r2302 := r2297(1 to 1);
    r2303 := r2297(2 to 2);
    r2304 := r2297(3 to 3);
    r2305 := r2297(4 to 4);
    r2306 := r2297(5 to 5);
    r2307 := r2297(6 to 6);
    r2308 := r2297(7 to 7);
    r2309 := r2297(8 to 8);
    r2310 := r2297(9 to 9);
    r2311 := r2297(10 to 10);
    r2312 := r2297(11 to 11);
    r2313 := r2297(12 to 12);
    r2314 := r2297(13 to 13);
    r2315 := r2297(14 to 14);
    r2316 := r2297(15 to 15);
    r2317 := r2297(16 to 16);
    r2318 := r2297(17 to 17);
    r2319 := r2297(18 to 18);
    r2320 := r2297(19 to 19);
    r2321 := r2297(20 to 20);
    r2322 := r2297(21 to 21);
    r2323 := r2297(22 to 22);
    r2324 := r2297(23 to 23);
    r2325 := r2297(24 to 24);
    r2326 := r2297(25 to 25);
    r2327 := r2297(26 to 26);
    r2328 := r2297(27 to 27);
    r2329 := r2297(28 to 28);
    r2330 := r2297(29 to 29);
    r2331 := r2297(30 to 30);
    r2332 := r2297(31 to 31);
    b2333 := true;
    b2334 := true;
    b2335 := true;
    b2336 := true;
    b2337 := true;
    b2338 := true;
    b2339 := true;
    b2340 := true;
    b2341 := true;
    b2342 := true;
    b2343 := true;
    b2344 := true;
    b2345 := true;
    b2346 := true;
    b2347 := true;
    b2348 := true;
    b2349 := true;
    b2350 := true;
    b2351 := true;
    b2352 := true;
    b2353 := true;
    b2354 := true;
    b2355 := true;
    b2356 := true;
    b2357 := true;
    b2358 := true;
    b2359 := true;
    b2360 := true;
    b2361 := true;
    b2362 := true;
    b2363 := true;
    b2364 := true;
    b2365 := (b2333 AND (b2334 AND (b2335 AND (b2336 AND (b2337 AND (b2338 AND (b2339 AND (b2340 AND (b2341 AND (b2342 AND (b2343 AND (b2344 AND (b2345 AND (b2346 AND (b2347 AND (b2348 AND (b2349 AND (b2350 AND (b2351 AND (b2352 AND (b2353 AND (b2354 AND (b2355 AND (b2356 AND (b2357 AND (b2358 AND (b2359 AND (b2360 AND (b2361 AND (b2362 AND (b2363 AND b2364)))))))))))))))))))))))))))))));
    if b2365 then
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      r2367 := (r2319 & r2320 & r2321 & r2322 & r2323 & r2324 & r2325 & r2326 & r2327 & r2328 & r2329 & r2330 & r2331 & r2332 & r2301 & r2302 & r2303 & r2304 & r2305 & r2306 & r2307 & r2308 & r2309 & r2310 & r2311 & r2312 & r2313 & r2314 & r2315 & r2316 & r2317 & r2318);
      r2299 := r2367;
    end if;
    return r2299;
  end rewire_rot18_2296;
  function rewire_rot13_2221(r2222 : std_logic_vector) return std_logic_vector
  is
    variable r2292 : std_logic_vector(0 to 31) := (others => '0');
    variable b2290 : boolean := false;
    variable b2289 : boolean := false;
    variable b2288 : boolean := false;
    variable b2287 : boolean := false;
    variable b2286 : boolean := false;
    variable b2285 : boolean := false;
    variable b2284 : boolean := false;
    variable b2283 : boolean := false;
    variable b2282 : boolean := false;
    variable b2281 : boolean := false;
    variable b2280 : boolean := false;
    variable b2279 : boolean := false;
    variable b2278 : boolean := false;
    variable b2277 : boolean := false;
    variable b2276 : boolean := false;
    variable b2275 : boolean := false;
    variable b2274 : boolean := false;
    variable b2273 : boolean := false;
    variable b2272 : boolean := false;
    variable b2271 : boolean := false;
    variable b2270 : boolean := false;
    variable b2269 : boolean := false;
    variable b2268 : boolean := false;
    variable b2267 : boolean := false;
    variable b2266 : boolean := false;
    variable b2265 : boolean := false;
    variable b2264 : boolean := false;
    variable b2263 : boolean := false;
    variable b2262 : boolean := false;
    variable b2261 : boolean := false;
    variable b2260 : boolean := false;
    variable b2259 : boolean := false;
    variable b2258 : boolean := false;
    variable r2257 : std_logic_vector(0 to 0) := (others => '0');
    variable r2256 : std_logic_vector(0 to 0) := (others => '0');
    variable r2255 : std_logic_vector(0 to 0) := (others => '0');
    variable r2254 : std_logic_vector(0 to 0) := (others => '0');
    variable r2253 : std_logic_vector(0 to 0) := (others => '0');
    variable r2252 : std_logic_vector(0 to 0) := (others => '0');
    variable r2251 : std_logic_vector(0 to 0) := (others => '0');
    variable r2250 : std_logic_vector(0 to 0) := (others => '0');
    variable r2249 : std_logic_vector(0 to 0) := (others => '0');
    variable r2248 : std_logic_vector(0 to 0) := (others => '0');
    variable r2247 : std_logic_vector(0 to 0) := (others => '0');
    variable r2246 : std_logic_vector(0 to 0) := (others => '0');
    variable r2245 : std_logic_vector(0 to 0) := (others => '0');
    variable r2244 : std_logic_vector(0 to 0) := (others => '0');
    variable r2243 : std_logic_vector(0 to 0) := (others => '0');
    variable r2242 : std_logic_vector(0 to 0) := (others => '0');
    variable r2241 : std_logic_vector(0 to 0) := (others => '0');
    variable r2240 : std_logic_vector(0 to 0) := (others => '0');
    variable r2239 : std_logic_vector(0 to 0) := (others => '0');
    variable r2238 : std_logic_vector(0 to 0) := (others => '0');
    variable r2237 : std_logic_vector(0 to 0) := (others => '0');
    variable r2236 : std_logic_vector(0 to 0) := (others => '0');
    variable r2235 : std_logic_vector(0 to 0) := (others => '0');
    variable r2234 : std_logic_vector(0 to 0) := (others => '0');
    variable r2233 : std_logic_vector(0 to 0) := (others => '0');
    variable r2232 : std_logic_vector(0 to 0) := (others => '0');
    variable r2231 : std_logic_vector(0 to 0) := (others => '0');
    variable r2230 : std_logic_vector(0 to 0) := (others => '0');
    variable r2229 : std_logic_vector(0 to 0) := (others => '0');
    variable r2228 : std_logic_vector(0 to 0) := (others => '0');
    variable r2227 : std_logic_vector(0 to 0) := (others => '0');
    variable r2226 : std_logic_vector(0 to 0) := (others => '0');
    variable b2225 : boolean := false;
    variable r2224 : std_logic_vector(0 to 31) := (others => '0');
  begin
    b2225 := true;
    r2226 := r2222(0 to 0);
    r2227 := r2222(1 to 1);
    r2228 := r2222(2 to 2);
    r2229 := r2222(3 to 3);
    r2230 := r2222(4 to 4);
    r2231 := r2222(5 to 5);
    r2232 := r2222(6 to 6);
    r2233 := r2222(7 to 7);
    r2234 := r2222(8 to 8);
    r2235 := r2222(9 to 9);
    r2236 := r2222(10 to 10);
    r2237 := r2222(11 to 11);
    r2238 := r2222(12 to 12);
    r2239 := r2222(13 to 13);
    r2240 := r2222(14 to 14);
    r2241 := r2222(15 to 15);
    r2242 := r2222(16 to 16);
    r2243 := r2222(17 to 17);
    r2244 := r2222(18 to 18);
    r2245 := r2222(19 to 19);
    r2246 := r2222(20 to 20);
    r2247 := r2222(21 to 21);
    r2248 := r2222(22 to 22);
    r2249 := r2222(23 to 23);
    r2250 := r2222(24 to 24);
    r2251 := r2222(25 to 25);
    r2252 := r2222(26 to 26);
    r2253 := r2222(27 to 27);
    r2254 := r2222(28 to 28);
    r2255 := r2222(29 to 29);
    r2256 := r2222(30 to 30);
    r2257 := r2222(31 to 31);
    b2258 := true;
    b2259 := true;
    b2260 := true;
    b2261 := true;
    b2262 := true;
    b2263 := true;
    b2264 := true;
    b2265 := true;
    b2266 := true;
    b2267 := true;
    b2268 := true;
    b2269 := true;
    b2270 := true;
    b2271 := true;
    b2272 := true;
    b2273 := true;
    b2274 := true;
    b2275 := true;
    b2276 := true;
    b2277 := true;
    b2278 := true;
    b2279 := true;
    b2280 := true;
    b2281 := true;
    b2282 := true;
    b2283 := true;
    b2284 := true;
    b2285 := true;
    b2286 := true;
    b2287 := true;
    b2288 := true;
    b2289 := true;
    b2290 := (b2258 AND (b2259 AND (b2260 AND (b2261 AND (b2262 AND (b2263 AND (b2264 AND (b2265 AND (b2266 AND (b2267 AND (b2268 AND (b2269 AND (b2270 AND (b2271 AND (b2272 AND (b2273 AND (b2274 AND (b2275 AND (b2276 AND (b2277 AND (b2278 AND (b2279 AND (b2280 AND (b2281 AND (b2282 AND (b2283 AND (b2284 AND (b2285 AND (b2286 AND (b2287 AND (b2288 AND b2289)))))))))))))))))))))))))))))));
    if b2290 then
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      r2292 := (r2239 & r2240 & r2241 & r2242 & r2243 & r2244 & r2245 & r2246 & r2247 & r2248 & r2249 & r2250 & r2251 & r2252 & r2253 & r2254 & r2255 & r2256 & r2257 & r2226 & r2227 & r2228 & r2229 & r2230 & r2231 & r2232 & r2233 & r2234 & r2235 & r2236 & r2237 & r2238);
      r2224 := r2292;
    end if;
    return r2224;
  end rewire_rot13_2221;
  function rewire_rot9_2146(r2147 : std_logic_vector) return std_logic_vector
  is
    variable r2217 : std_logic_vector(0 to 31) := (others => '0');
    variable b2215 : boolean := false;
    variable b2214 : boolean := false;
    variable b2213 : boolean := false;
    variable b2212 : boolean := false;
    variable b2211 : boolean := false;
    variable b2210 : boolean := false;
    variable b2209 : boolean := false;
    variable b2208 : boolean := false;
    variable b2207 : boolean := false;
    variable b2206 : boolean := false;
    variable b2205 : boolean := false;
    variable b2204 : boolean := false;
    variable b2203 : boolean := false;
    variable b2202 : boolean := false;
    variable b2201 : boolean := false;
    variable b2200 : boolean := false;
    variable b2199 : boolean := false;
    variable b2198 : boolean := false;
    variable b2197 : boolean := false;
    variable b2196 : boolean := false;
    variable b2195 : boolean := false;
    variable b2194 : boolean := false;
    variable b2193 : boolean := false;
    variable b2192 : boolean := false;
    variable b2191 : boolean := false;
    variable b2190 : boolean := false;
    variable b2189 : boolean := false;
    variable b2188 : boolean := false;
    variable b2187 : boolean := false;
    variable b2186 : boolean := false;
    variable b2185 : boolean := false;
    variable b2184 : boolean := false;
    variable b2183 : boolean := false;
    variable r2182 : std_logic_vector(0 to 0) := (others => '0');
    variable r2181 : std_logic_vector(0 to 0) := (others => '0');
    variable r2180 : std_logic_vector(0 to 0) := (others => '0');
    variable r2179 : std_logic_vector(0 to 0) := (others => '0');
    variable r2178 : std_logic_vector(0 to 0) := (others => '0');
    variable r2177 : std_logic_vector(0 to 0) := (others => '0');
    variable r2176 : std_logic_vector(0 to 0) := (others => '0');
    variable r2175 : std_logic_vector(0 to 0) := (others => '0');
    variable r2174 : std_logic_vector(0 to 0) := (others => '0');
    variable r2173 : std_logic_vector(0 to 0) := (others => '0');
    variable r2172 : std_logic_vector(0 to 0) := (others => '0');
    variable r2171 : std_logic_vector(0 to 0) := (others => '0');
    variable r2170 : std_logic_vector(0 to 0) := (others => '0');
    variable r2169 : std_logic_vector(0 to 0) := (others => '0');
    variable r2168 : std_logic_vector(0 to 0) := (others => '0');
    variable r2167 : std_logic_vector(0 to 0) := (others => '0');
    variable r2166 : std_logic_vector(0 to 0) := (others => '0');
    variable r2165 : std_logic_vector(0 to 0) := (others => '0');
    variable r2164 : std_logic_vector(0 to 0) := (others => '0');
    variable r2163 : std_logic_vector(0 to 0) := (others => '0');
    variable r2162 : std_logic_vector(0 to 0) := (others => '0');
    variable r2161 : std_logic_vector(0 to 0) := (others => '0');
    variable r2160 : std_logic_vector(0 to 0) := (others => '0');
    variable r2159 : std_logic_vector(0 to 0) := (others => '0');
    variable r2158 : std_logic_vector(0 to 0) := (others => '0');
    variable r2157 : std_logic_vector(0 to 0) := (others => '0');
    variable r2156 : std_logic_vector(0 to 0) := (others => '0');
    variable r2155 : std_logic_vector(0 to 0) := (others => '0');
    variable r2154 : std_logic_vector(0 to 0) := (others => '0');
    variable r2153 : std_logic_vector(0 to 0) := (others => '0');
    variable r2152 : std_logic_vector(0 to 0) := (others => '0');
    variable r2151 : std_logic_vector(0 to 0) := (others => '0');
    variable b2150 : boolean := false;
    variable r2149 : std_logic_vector(0 to 31) := (others => '0');
  begin
    b2150 := true;
    r2151 := r2147(0 to 0);
    r2152 := r2147(1 to 1);
    r2153 := r2147(2 to 2);
    r2154 := r2147(3 to 3);
    r2155 := r2147(4 to 4);
    r2156 := r2147(5 to 5);
    r2157 := r2147(6 to 6);
    r2158 := r2147(7 to 7);
    r2159 := r2147(8 to 8);
    r2160 := r2147(9 to 9);
    r2161 := r2147(10 to 10);
    r2162 := r2147(11 to 11);
    r2163 := r2147(12 to 12);
    r2164 := r2147(13 to 13);
    r2165 := r2147(14 to 14);
    r2166 := r2147(15 to 15);
    r2167 := r2147(16 to 16);
    r2168 := r2147(17 to 17);
    r2169 := r2147(18 to 18);
    r2170 := r2147(19 to 19);
    r2171 := r2147(20 to 20);
    r2172 := r2147(21 to 21);
    r2173 := r2147(22 to 22);
    r2174 := r2147(23 to 23);
    r2175 := r2147(24 to 24);
    r2176 := r2147(25 to 25);
    r2177 := r2147(26 to 26);
    r2178 := r2147(27 to 27);
    r2179 := r2147(28 to 28);
    r2180 := r2147(29 to 29);
    r2181 := r2147(30 to 30);
    r2182 := r2147(31 to 31);
    b2183 := true;
    b2184 := true;
    b2185 := true;
    b2186 := true;
    b2187 := true;
    b2188 := true;
    b2189 := true;
    b2190 := true;
    b2191 := true;
    b2192 := true;
    b2193 := true;
    b2194 := true;
    b2195 := true;
    b2196 := true;
    b2197 := true;
    b2198 := true;
    b2199 := true;
    b2200 := true;
    b2201 := true;
    b2202 := true;
    b2203 := true;
    b2204 := true;
    b2205 := true;
    b2206 := true;
    b2207 := true;
    b2208 := true;
    b2209 := true;
    b2210 := true;
    b2211 := true;
    b2212 := true;
    b2213 := true;
    b2214 := true;
    b2215 := (b2183 AND (b2184 AND (b2185 AND (b2186 AND (b2187 AND (b2188 AND (b2189 AND (b2190 AND (b2191 AND (b2192 AND (b2193 AND (b2194 AND (b2195 AND (b2196 AND (b2197 AND (b2198 AND (b2199 AND (b2200 AND (b2201 AND (b2202 AND (b2203 AND (b2204 AND (b2205 AND (b2206 AND (b2207 AND (b2208 AND (b2209 AND (b2210 AND (b2211 AND (b2212 AND (b2213 AND b2214)))))))))))))))))))))))))))))));
    if b2215 then
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      r2217 := (r2160 & r2161 & r2162 & r2163 & r2164 & r2165 & r2166 & r2167 & r2168 & r2169 & r2170 & r2171 & r2172 & r2173 & r2174 & r2175 & r2176 & r2177 & r2178 & r2179 & r2180 & r2181 & r2182 & r2151 & r2152 & r2153 & r2154 & r2155 & r2156 & r2157 & r2158 & r2159);
      r2149 := r2217;
    end if;
    return r2149;
  end rewire_rot9_2146;
  function rewire_rot7_2071(r2072 : std_logic_vector) return std_logic_vector
  is
    variable r2142 : std_logic_vector(0 to 31) := (others => '0');
    variable b2140 : boolean := false;
    variable b2139 : boolean := false;
    variable b2138 : boolean := false;
    variable b2137 : boolean := false;
    variable b2136 : boolean := false;
    variable b2135 : boolean := false;
    variable b2134 : boolean := false;
    variable b2133 : boolean := false;
    variable b2132 : boolean := false;
    variable b2131 : boolean := false;
    variable b2130 : boolean := false;
    variable b2129 : boolean := false;
    variable b2128 : boolean := false;
    variable b2127 : boolean := false;
    variable b2126 : boolean := false;
    variable b2125 : boolean := false;
    variable b2124 : boolean := false;
    variable b2123 : boolean := false;
    variable b2122 : boolean := false;
    variable b2121 : boolean := false;
    variable b2120 : boolean := false;
    variable b2119 : boolean := false;
    variable b2118 : boolean := false;
    variable b2117 : boolean := false;
    variable b2116 : boolean := false;
    variable b2115 : boolean := false;
    variable b2114 : boolean := false;
    variable b2113 : boolean := false;
    variable b2112 : boolean := false;
    variable b2111 : boolean := false;
    variable b2110 : boolean := false;
    variable b2109 : boolean := false;
    variable b2108 : boolean := false;
    variable r2107 : std_logic_vector(0 to 0) := (others => '0');
    variable r2106 : std_logic_vector(0 to 0) := (others => '0');
    variable r2105 : std_logic_vector(0 to 0) := (others => '0');
    variable r2104 : std_logic_vector(0 to 0) := (others => '0');
    variable r2103 : std_logic_vector(0 to 0) := (others => '0');
    variable r2102 : std_logic_vector(0 to 0) := (others => '0');
    variable r2101 : std_logic_vector(0 to 0) := (others => '0');
    variable r2100 : std_logic_vector(0 to 0) := (others => '0');
    variable r2099 : std_logic_vector(0 to 0) := (others => '0');
    variable r2098 : std_logic_vector(0 to 0) := (others => '0');
    variable r2097 : std_logic_vector(0 to 0) := (others => '0');
    variable r2096 : std_logic_vector(0 to 0) := (others => '0');
    variable r2095 : std_logic_vector(0 to 0) := (others => '0');
    variable r2094 : std_logic_vector(0 to 0) := (others => '0');
    variable r2093 : std_logic_vector(0 to 0) := (others => '0');
    variable r2092 : std_logic_vector(0 to 0) := (others => '0');
    variable r2091 : std_logic_vector(0 to 0) := (others => '0');
    variable r2090 : std_logic_vector(0 to 0) := (others => '0');
    variable r2089 : std_logic_vector(0 to 0) := (others => '0');
    variable r2088 : std_logic_vector(0 to 0) := (others => '0');
    variable r2087 : std_logic_vector(0 to 0) := (others => '0');
    variable r2086 : std_logic_vector(0 to 0) := (others => '0');
    variable r2085 : std_logic_vector(0 to 0) := (others => '0');
    variable r2084 : std_logic_vector(0 to 0) := (others => '0');
    variable r2083 : std_logic_vector(0 to 0) := (others => '0');
    variable r2082 : std_logic_vector(0 to 0) := (others => '0');
    variable r2081 : std_logic_vector(0 to 0) := (others => '0');
    variable r2080 : std_logic_vector(0 to 0) := (others => '0');
    variable r2079 : std_logic_vector(0 to 0) := (others => '0');
    variable r2078 : std_logic_vector(0 to 0) := (others => '0');
    variable r2077 : std_logic_vector(0 to 0) := (others => '0');
    variable r2076 : std_logic_vector(0 to 0) := (others => '0');
    variable b2075 : boolean := false;
    variable r2074 : std_logic_vector(0 to 31) := (others => '0');
  begin
    b2075 := true;
    r2076 := r2072(0 to 0);
    r2077 := r2072(1 to 1);
    r2078 := r2072(2 to 2);
    r2079 := r2072(3 to 3);
    r2080 := r2072(4 to 4);
    r2081 := r2072(5 to 5);
    r2082 := r2072(6 to 6);
    r2083 := r2072(7 to 7);
    r2084 := r2072(8 to 8);
    r2085 := r2072(9 to 9);
    r2086 := r2072(10 to 10);
    r2087 := r2072(11 to 11);
    r2088 := r2072(12 to 12);
    r2089 := r2072(13 to 13);
    r2090 := r2072(14 to 14);
    r2091 := r2072(15 to 15);
    r2092 := r2072(16 to 16);
    r2093 := r2072(17 to 17);
    r2094 := r2072(18 to 18);
    r2095 := r2072(19 to 19);
    r2096 := r2072(20 to 20);
    r2097 := r2072(21 to 21);
    r2098 := r2072(22 to 22);
    r2099 := r2072(23 to 23);
    r2100 := r2072(24 to 24);
    r2101 := r2072(25 to 25);
    r2102 := r2072(26 to 26);
    r2103 := r2072(27 to 27);
    r2104 := r2072(28 to 28);
    r2105 := r2072(29 to 29);
    r2106 := r2072(30 to 30);
    r2107 := r2072(31 to 31);
    b2108 := true;
    b2109 := true;
    b2110 := true;
    b2111 := true;
    b2112 := true;
    b2113 := true;
    b2114 := true;
    b2115 := true;
    b2116 := true;
    b2117 := true;
    b2118 := true;
    b2119 := true;
    b2120 := true;
    b2121 := true;
    b2122 := true;
    b2123 := true;
    b2124 := true;
    b2125 := true;
    b2126 := true;
    b2127 := true;
    b2128 := true;
    b2129 := true;
    b2130 := true;
    b2131 := true;
    b2132 := true;
    b2133 := true;
    b2134 := true;
    b2135 := true;
    b2136 := true;
    b2137 := true;
    b2138 := true;
    b2139 := true;
    b2140 := (b2108 AND (b2109 AND (b2110 AND (b2111 AND (b2112 AND (b2113 AND (b2114 AND (b2115 AND (b2116 AND (b2117 AND (b2118 AND (b2119 AND (b2120 AND (b2121 AND (b2122 AND (b2123 AND (b2124 AND (b2125 AND (b2126 AND (b2127 AND (b2128 AND (b2129 AND (b2130 AND (b2131 AND (b2132 AND (b2133 AND (b2134 AND (b2135 AND (b2136 AND (b2137 AND (b2138 AND b2139)))))))))))))))))))))))))))))));
    if b2140 then
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      r2142 := (r2083 & r2084 & r2085 & r2086 & r2087 & r2088 & r2089 & r2090 & r2091 & r2092 & r2093 & r2094 & r2095 & r2096 & r2097 & r2098 & r2099 & r2100 & r2101 & r2102 & r2103 & r2104 & r2105 & r2106 & r2107 & r2076 & r2077 & r2078 & r2079 & r2080 & r2081 & r2082);
      r2074 := r2142;
    end if;
    return r2074;
  end rewire_rot7_2071;
  function rewire_expwords_1661(r1662 : std_logic_vector) return std_logic_vector
  is
    variable r1977 : std_logic_vector(0 to 511) := (others => '0');
    variable b1975 : boolean := false;
    variable b1974 : boolean := false;
    variable b1973 : boolean := false;
    variable b1972 : boolean := false;
    variable b1971 : boolean := false;
    variable b1970 : boolean := false;
    variable r1969 : std_logic_vector(0 to 7) := (others => '0');
    variable r1968 : std_logic_vector(0 to 7) := (others => '0');
    variable r1967 : std_logic_vector(0 to 7) := (others => '0');
    variable r1966 : std_logic_vector(0 to 7) := (others => '0');
    variable b1965 : boolean := false;
    variable b1964 : boolean := false;
    variable b1963 : boolean := false;
    variable b1962 : boolean := false;
    variable b1961 : boolean := false;
    variable b1960 : boolean := false;
    variable r1959 : std_logic_vector(0 to 7) := (others => '0');
    variable r1958 : std_logic_vector(0 to 7) := (others => '0');
    variable r1957 : std_logic_vector(0 to 7) := (others => '0');
    variable r1956 : std_logic_vector(0 to 7) := (others => '0');
    variable b1955 : boolean := false;
    variable b1954 : boolean := false;
    variable b1953 : boolean := false;
    variable b1952 : boolean := false;
    variable b1951 : boolean := false;
    variable b1950 : boolean := false;
    variable r1949 : std_logic_vector(0 to 7) := (others => '0');
    variable r1948 : std_logic_vector(0 to 7) := (others => '0');
    variable r1947 : std_logic_vector(0 to 7) := (others => '0');
    variable r1946 : std_logic_vector(0 to 7) := (others => '0');
    variable b1945 : boolean := false;
    variable b1944 : boolean := false;
    variable b1943 : boolean := false;
    variable b1942 : boolean := false;
    variable b1941 : boolean := false;
    variable b1940 : boolean := false;
    variable r1939 : std_logic_vector(0 to 7) := (others => '0');
    variable r1938 : std_logic_vector(0 to 7) := (others => '0');
    variable r1937 : std_logic_vector(0 to 7) := (others => '0');
    variable r1936 : std_logic_vector(0 to 7) := (others => '0');
    variable b1935 : boolean := false;
    variable b1934 : boolean := false;
    variable b1933 : boolean := false;
    variable b1932 : boolean := false;
    variable b1931 : boolean := false;
    variable b1930 : boolean := false;
    variable r1929 : std_logic_vector(0 to 7) := (others => '0');
    variable r1928 : std_logic_vector(0 to 7) := (others => '0');
    variable r1927 : std_logic_vector(0 to 7) := (others => '0');
    variable r1926 : std_logic_vector(0 to 7) := (others => '0');
    variable b1925 : boolean := false;
    variable b1924 : boolean := false;
    variable b1923 : boolean := false;
    variable b1922 : boolean := false;
    variable b1921 : boolean := false;
    variable b1920 : boolean := false;
    variable r1919 : std_logic_vector(0 to 7) := (others => '0');
    variable r1918 : std_logic_vector(0 to 7) := (others => '0');
    variable r1917 : std_logic_vector(0 to 7) := (others => '0');
    variable r1916 : std_logic_vector(0 to 7) := (others => '0');
    variable b1915 : boolean := false;
    variable b1914 : boolean := false;
    variable b1913 : boolean := false;
    variable b1912 : boolean := false;
    variable b1911 : boolean := false;
    variable b1910 : boolean := false;
    variable r1909 : std_logic_vector(0 to 7) := (others => '0');
    variable r1908 : std_logic_vector(0 to 7) := (others => '0');
    variable r1907 : std_logic_vector(0 to 7) := (others => '0');
    variable r1906 : std_logic_vector(0 to 7) := (others => '0');
    variable b1905 : boolean := false;
    variable b1904 : boolean := false;
    variable b1903 : boolean := false;
    variable b1902 : boolean := false;
    variable b1901 : boolean := false;
    variable b1900 : boolean := false;
    variable r1899 : std_logic_vector(0 to 7) := (others => '0');
    variable r1898 : std_logic_vector(0 to 7) := (others => '0');
    variable r1897 : std_logic_vector(0 to 7) := (others => '0');
    variable r1896 : std_logic_vector(0 to 7) := (others => '0');
    variable b1895 : boolean := false;
    variable b1894 : boolean := false;
    variable b1893 : boolean := false;
    variable b1892 : boolean := false;
    variable b1891 : boolean := false;
    variable b1890 : boolean := false;
    variable r1889 : std_logic_vector(0 to 7) := (others => '0');
    variable r1888 : std_logic_vector(0 to 7) := (others => '0');
    variable r1887 : std_logic_vector(0 to 7) := (others => '0');
    variable r1886 : std_logic_vector(0 to 7) := (others => '0');
    variable b1885 : boolean := false;
    variable b1884 : boolean := false;
    variable b1883 : boolean := false;
    variable b1882 : boolean := false;
    variable b1881 : boolean := false;
    variable b1880 : boolean := false;
    variable r1879 : std_logic_vector(0 to 7) := (others => '0');
    variable r1878 : std_logic_vector(0 to 7) := (others => '0');
    variable r1877 : std_logic_vector(0 to 7) := (others => '0');
    variable r1876 : std_logic_vector(0 to 7) := (others => '0');
    variable b1875 : boolean := false;
    variable b1874 : boolean := false;
    variable b1873 : boolean := false;
    variable b1872 : boolean := false;
    variable b1871 : boolean := false;
    variable b1870 : boolean := false;
    variable r1869 : std_logic_vector(0 to 7) := (others => '0');
    variable r1868 : std_logic_vector(0 to 7) := (others => '0');
    variable r1867 : std_logic_vector(0 to 7) := (others => '0');
    variable r1866 : std_logic_vector(0 to 7) := (others => '0');
    variable b1865 : boolean := false;
    variable b1864 : boolean := false;
    variable b1863 : boolean := false;
    variable b1862 : boolean := false;
    variable b1861 : boolean := false;
    variable b1860 : boolean := false;
    variable r1859 : std_logic_vector(0 to 7) := (others => '0');
    variable r1858 : std_logic_vector(0 to 7) := (others => '0');
    variable r1857 : std_logic_vector(0 to 7) := (others => '0');
    variable r1856 : std_logic_vector(0 to 7) := (others => '0');
    variable b1855 : boolean := false;
    variable b1854 : boolean := false;
    variable b1853 : boolean := false;
    variable b1852 : boolean := false;
    variable b1851 : boolean := false;
    variable b1850 : boolean := false;
    variable r1849 : std_logic_vector(0 to 7) := (others => '0');
    variable r1848 : std_logic_vector(0 to 7) := (others => '0');
    variable r1847 : std_logic_vector(0 to 7) := (others => '0');
    variable r1846 : std_logic_vector(0 to 7) := (others => '0');
    variable b1845 : boolean := false;
    variable b1844 : boolean := false;
    variable b1843 : boolean := false;
    variable b1842 : boolean := false;
    variable b1841 : boolean := false;
    variable b1840 : boolean := false;
    variable r1839 : std_logic_vector(0 to 7) := (others => '0');
    variable r1838 : std_logic_vector(0 to 7) := (others => '0');
    variable r1837 : std_logic_vector(0 to 7) := (others => '0');
    variable r1836 : std_logic_vector(0 to 7) := (others => '0');
    variable b1835 : boolean := false;
    variable b1834 : boolean := false;
    variable b1833 : boolean := false;
    variable b1832 : boolean := false;
    variable b1831 : boolean := false;
    variable b1830 : boolean := false;
    variable r1829 : std_logic_vector(0 to 7) := (others => '0');
    variable r1828 : std_logic_vector(0 to 7) := (others => '0');
    variable r1827 : std_logic_vector(0 to 7) := (others => '0');
    variable r1826 : std_logic_vector(0 to 7) := (others => '0');
    variable b1825 : boolean := false;
    variable b1824 : boolean := false;
    variable b1823 : boolean := false;
    variable b1822 : boolean := false;
    variable b1821 : boolean := false;
    variable b1820 : boolean := false;
    variable r1819 : std_logic_vector(0 to 7) := (others => '0');
    variable r1818 : std_logic_vector(0 to 7) := (others => '0');
    variable r1817 : std_logic_vector(0 to 7) := (others => '0');
    variable r1816 : std_logic_vector(0 to 7) := (others => '0');
    variable b1815 : boolean := false;
    variable r1814 : std_logic_vector(0 to 31) := (others => '0');
    variable r1813 : std_logic_vector(0 to 31) := (others => '0');
    variable r1812 : std_logic_vector(0 to 31) := (others => '0');
    variable r1811 : std_logic_vector(0 to 31) := (others => '0');
    variable r1810 : std_logic_vector(0 to 31) := (others => '0');
    variable r1809 : std_logic_vector(0 to 31) := (others => '0');
    variable r1808 : std_logic_vector(0 to 31) := (others => '0');
    variable r1807 : std_logic_vector(0 to 31) := (others => '0');
    variable r1806 : std_logic_vector(0 to 31) := (others => '0');
    variable r1805 : std_logic_vector(0 to 31) := (others => '0');
    variable r1804 : std_logic_vector(0 to 31) := (others => '0');
    variable r1803 : std_logic_vector(0 to 31) := (others => '0');
    variable r1802 : std_logic_vector(0 to 31) := (others => '0');
    variable r1801 : std_logic_vector(0 to 31) := (others => '0');
    variable r1800 : std_logic_vector(0 to 31) := (others => '0');
    variable r1799 : std_logic_vector(0 to 31) := (others => '0');
    variable b1798 : boolean := false;
    variable r1797 : std_logic_vector(0 to 511) := (others => '0');
    variable r1796 : std_logic_vector(0 to 511) := (others => '0');
    variable r1794 : std_logic_vector(0 to 31) := (others => '0');
    variable r1793 : std_logic_vector(0 to 31) := (others => '0');
    variable r1792 : std_logic_vector(0 to 31) := (others => '0');
    variable r1791 : std_logic_vector(0 to 31) := (others => '0');
    variable r1790 : std_logic_vector(0 to 31) := (others => '0');
    variable r1789 : std_logic_vector(0 to 31) := (others => '0');
    variable r1788 : std_logic_vector(0 to 31) := (others => '0');
    variable r1787 : std_logic_vector(0 to 31) := (others => '0');
    variable r1786 : std_logic_vector(0 to 31) := (others => '0');
    variable r1785 : std_logic_vector(0 to 31) := (others => '0');
    variable r1784 : std_logic_vector(0 to 31) := (others => '0');
    variable r1783 : std_logic_vector(0 to 31) := (others => '0');
    variable r1782 : std_logic_vector(0 to 31) := (others => '0');
    variable r1781 : std_logic_vector(0 to 31) := (others => '0');
    variable r1780 : std_logic_vector(0 to 31) := (others => '0');
    variable r1779 : std_logic_vector(0 to 31) := (others => '0');
    variable r1701 : std_logic_vector(0 to 31) := (others => '0');
    variable r1700 : std_logic_vector(0 to 31) := (others => '0');
    variable b1698 : boolean := false;
    variable b1697 : boolean := false;
    variable b1696 : boolean := false;
    variable b1695 : boolean := false;
    variable b1694 : boolean := false;
    variable b1693 : boolean := false;
    variable b1692 : boolean := false;
    variable b1691 : boolean := false;
    variable b1690 : boolean := false;
    variable b1689 : boolean := false;
    variable b1688 : boolean := false;
    variable b1687 : boolean := false;
    variable b1686 : boolean := false;
    variable b1685 : boolean := false;
    variable b1684 : boolean := false;
    variable b1683 : boolean := false;
    variable b1682 : boolean := false;
    variable r1681 : std_logic_vector(0 to 31) := (others => '0');
    variable r1680 : std_logic_vector(0 to 31) := (others => '0');
    variable r1679 : std_logic_vector(0 to 31) := (others => '0');
    variable r1678 : std_logic_vector(0 to 31) := (others => '0');
    variable r1677 : std_logic_vector(0 to 31) := (others => '0');
    variable r1676 : std_logic_vector(0 to 31) := (others => '0');
    variable r1675 : std_logic_vector(0 to 31) := (others => '0');
    variable r1674 : std_logic_vector(0 to 31) := (others => '0');
    variable r1673 : std_logic_vector(0 to 31) := (others => '0');
    variable r1672 : std_logic_vector(0 to 31) := (others => '0');
    variable r1671 : std_logic_vector(0 to 31) := (others => '0');
    variable r1670 : std_logic_vector(0 to 31) := (others => '0');
    variable r1669 : std_logic_vector(0 to 31) := (others => '0');
    variable r1668 : std_logic_vector(0 to 31) := (others => '0');
    variable r1667 : std_logic_vector(0 to 31) := (others => '0');
    variable r1666 : std_logic_vector(0 to 31) := (others => '0');
    variable b1665 : boolean := false;
    variable r1664 : std_logic_vector(0 to 511) := (others => '0');
  begin
    b1665 := true;
    r1666 := r1662(0 to 31);
    r1667 := r1662(32 to 63);
    r1668 := r1662(64 to 95);
    r1669 := r1662(96 to 127);
    r1670 := r1662(128 to 159);
    r1671 := r1662(160 to 191);
    r1672 := r1662(192 to 223);
    r1673 := r1662(224 to 255);
    r1674 := r1662(256 to 287);
    r1675 := r1662(288 to 319);
    r1676 := r1662(320 to 351);
    r1677 := r1662(352 to 383);
    r1678 := r1662(384 to 415);
    r1679 := r1662(416 to 447);
    r1680 := r1662(448 to 479);
    r1681 := r1662(480 to 511);
    b1682 := true;
    b1683 := true;
    b1684 := true;
    b1685 := true;
    b1686 := true;
    b1687 := true;
    b1688 := true;
    b1689 := true;
    b1690 := true;
    b1691 := true;
    b1692 := true;
    b1693 := true;
    b1694 := true;
    b1695 := true;
    b1696 := true;
    b1697 := true;
    b1698 := (b1682 AND (b1683 AND (b1684 AND (b1685 AND (b1686 AND (b1687 AND (b1688 AND (b1689 AND (b1690 AND (b1691 AND (b1692 AND (b1693 AND (b1694 AND (b1695 AND (b1696 AND b1697)))))))))))))));
    if b1698 then
      null;
      r1779 := rewire_littleendianp_1699(r1666);
      null;
      r1780 := rewire_littleendianp_1699(r1667);
      null;
      r1781 := rewire_littleendianp_1699(r1668);
      null;
      r1782 := rewire_littleendianp_1699(r1669);
      null;
      r1783 := rewire_littleendianp_1699(r1670);
      null;
      r1784 := rewire_littleendianp_1699(r1671);
      null;
      r1785 := rewire_littleendianp_1699(r1672);
      null;
      r1786 := rewire_littleendianp_1699(r1673);
      null;
      r1787 := rewire_littleendianp_1699(r1674);
      null;
      r1788 := rewire_littleendianp_1699(r1675);
      null;
      r1789 := rewire_littleendianp_1699(r1676);
      null;
      r1790 := rewire_littleendianp_1699(r1677);
      null;
      r1791 := rewire_littleendianp_1699(r1678);
      null;
      r1792 := rewire_littleendianp_1699(r1679);
      null;
      r1793 := rewire_littleendianp_1699(r1680);
      null;
      r1794 := rewire_littleendianp_1699(r1681);
      b1798 := true;
      r1799 := r1796(0 to 31);
      r1800 := r1796(32 to 63);
      r1801 := r1796(64 to 95);
      r1802 := r1796(96 to 127);
      r1803 := r1796(128 to 159);
      r1804 := r1796(160 to 191);
      r1805 := r1796(192 to 223);
      r1806 := r1796(224 to 255);
      r1807 := r1796(256 to 287);
      r1808 := r1796(288 to 319);
      r1809 := r1796(320 to 351);
      r1810 := r1796(352 to 383);
      r1811 := r1796(384 to 415);
      r1812 := r1796(416 to 447);
      r1813 := r1796(448 to 479);
      r1814 := r1796(480 to 511);
      b1815 := true;
      r1816 := r1799(0 to 7);
      r1817 := r1799(8 to 15);
      r1818 := r1799(16 to 23);
      r1819 := r1799(24 to 31);
      b1820 := true;
      b1821 := true;
      b1822 := true;
      b1823 := true;
      b1824 := (b1820 AND (b1821 AND (b1822 AND b1823)));
      b1825 := true;
      r1826 := r1800(0 to 7);
      r1827 := r1800(8 to 15);
      r1828 := r1800(16 to 23);
      r1829 := r1800(24 to 31);
      b1830 := true;
      b1831 := true;
      b1832 := true;
      b1833 := true;
      b1834 := (b1830 AND (b1831 AND (b1832 AND b1833)));
      b1835 := true;
      r1836 := r1801(0 to 7);
      r1837 := r1801(8 to 15);
      r1838 := r1801(16 to 23);
      r1839 := r1801(24 to 31);
      b1840 := true;
      b1841 := true;
      b1842 := true;
      b1843 := true;
      b1844 := (b1840 AND (b1841 AND (b1842 AND b1843)));
      b1845 := true;
      r1846 := r1802(0 to 7);
      r1847 := r1802(8 to 15);
      r1848 := r1802(16 to 23);
      r1849 := r1802(24 to 31);
      b1850 := true;
      b1851 := true;
      b1852 := true;
      b1853 := true;
      b1854 := (b1850 AND (b1851 AND (b1852 AND b1853)));
      b1855 := true;
      r1856 := r1803(0 to 7);
      r1857 := r1803(8 to 15);
      r1858 := r1803(16 to 23);
      r1859 := r1803(24 to 31);
      b1860 := true;
      b1861 := true;
      b1862 := true;
      b1863 := true;
      b1864 := (b1860 AND (b1861 AND (b1862 AND b1863)));
      b1865 := true;
      r1866 := r1804(0 to 7);
      r1867 := r1804(8 to 15);
      r1868 := r1804(16 to 23);
      r1869 := r1804(24 to 31);
      b1870 := true;
      b1871 := true;
      b1872 := true;
      b1873 := true;
      b1874 := (b1870 AND (b1871 AND (b1872 AND b1873)));
      b1875 := true;
      r1876 := r1805(0 to 7);
      r1877 := r1805(8 to 15);
      r1878 := r1805(16 to 23);
      r1879 := r1805(24 to 31);
      b1880 := true;
      b1881 := true;
      b1882 := true;
      b1883 := true;
      b1884 := (b1880 AND (b1881 AND (b1882 AND b1883)));
      b1885 := true;
      r1886 := r1806(0 to 7);
      r1887 := r1806(8 to 15);
      r1888 := r1806(16 to 23);
      r1889 := r1806(24 to 31);
      b1890 := true;
      b1891 := true;
      b1892 := true;
      b1893 := true;
      b1894 := (b1890 AND (b1891 AND (b1892 AND b1893)));
      b1895 := true;
      r1896 := r1807(0 to 7);
      r1897 := r1807(8 to 15);
      r1898 := r1807(16 to 23);
      r1899 := r1807(24 to 31);
      b1900 := true;
      b1901 := true;
      b1902 := true;
      b1903 := true;
      b1904 := (b1900 AND (b1901 AND (b1902 AND b1903)));
      b1905 := true;
      r1906 := r1808(0 to 7);
      r1907 := r1808(8 to 15);
      r1908 := r1808(16 to 23);
      r1909 := r1808(24 to 31);
      b1910 := true;
      b1911 := true;
      b1912 := true;
      b1913 := true;
      b1914 := (b1910 AND (b1911 AND (b1912 AND b1913)));
      b1915 := true;
      r1916 := r1809(0 to 7);
      r1917 := r1809(8 to 15);
      r1918 := r1809(16 to 23);
      r1919 := r1809(24 to 31);
      b1920 := true;
      b1921 := true;
      b1922 := true;
      b1923 := true;
      b1924 := (b1920 AND (b1921 AND (b1922 AND b1923)));
      b1925 := true;
      r1926 := r1810(0 to 7);
      r1927 := r1810(8 to 15);
      r1928 := r1810(16 to 23);
      r1929 := r1810(24 to 31);
      b1930 := true;
      b1931 := true;
      b1932 := true;
      b1933 := true;
      b1934 := (b1930 AND (b1931 AND (b1932 AND b1933)));
      b1935 := true;
      r1936 := r1811(0 to 7);
      r1937 := r1811(8 to 15);
      r1938 := r1811(16 to 23);
      r1939 := r1811(24 to 31);
      b1940 := true;
      b1941 := true;
      b1942 := true;
      b1943 := true;
      b1944 := (b1940 AND (b1941 AND (b1942 AND b1943)));
      b1945 := true;
      r1946 := r1812(0 to 7);
      r1947 := r1812(8 to 15);
      r1948 := r1812(16 to 23);
      r1949 := r1812(24 to 31);
      b1950 := true;
      b1951 := true;
      b1952 := true;
      b1953 := true;
      b1954 := (b1950 AND (b1951 AND (b1952 AND b1953)));
      b1955 := true;
      r1956 := r1813(0 to 7);
      r1957 := r1813(8 to 15);
      r1958 := r1813(16 to 23);
      r1959 := r1813(24 to 31);
      b1960 := true;
      b1961 := true;
      b1962 := true;
      b1963 := true;
      b1964 := (b1960 AND (b1961 AND (b1962 AND b1963)));
      b1965 := true;
      r1966 := r1814(0 to 7);
      r1967 := r1814(8 to 15);
      r1968 := r1814(16 to 23);
      r1969 := r1814(24 to 31);
      b1970 := true;
      b1971 := true;
      b1972 := true;
      b1973 := true;
      b1974 := (b1970 AND (b1971 AND (b1972 AND b1973)));
      b1975 := (b1824 AND (b1834 AND (b1844 AND (b1854 AND (b1864 AND (b1874 AND (b1884 AND (b1894 AND (b1904 AND (b1914 AND (b1924 AND (b1934 AND (b1944 AND (b1954 AND (b1964 AND b1974)))))))))))))));
      if b1975 then
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        r1977 := (r1816 & r1817 & r1818 & r1819 & r1826 & r1827 & r1828 & r1829 & r1836 & r1837 & r1838 & r1839 & r1846 & r1847 & r1848 & r1849 & r1856 & r1857 & r1858 & r1859 & r1866 & r1867 & r1868 & r1869 & r1876 & r1877 & r1878 & r1879 & r1886 & r1887 & r1888 & r1889 & r1896 & r1897 & r1898 & r1899 & r1906 & r1907 & r1908 & r1909 & r1916 & r1917 & r1918 & r1919 & r1926 & r1927 & r1928 & r1929 & r1936 & r1937 & r1938 & r1939 & r1946 & r1947 & r1948 & r1949 & r1956 & r1957 & r1958 & r1959 & r1966 & r1967 & r1968 & r1969);
        r1797 := r1977;
      end if;
      r1664 := r1797;
    end if;
    return r1664;
  end rewire_expwords_1661;
  function rewire_littleendianp_1699(r1700 : std_logic_vector) return std_logic_vector
  is
    variable r1778 : std_logic_vector(0 to 31) := (others => '0');
    variable r1777 : std_logic_vector(0 to 7) := (others => '0');
    variable r1775 : std_logic_vector(0 to 7) := (others => '0');
    variable r1773 : std_logic_vector(0 to 7) := (others => '0');
    variable r1771 : std_logic_vector(0 to 7) := (others => '0');
    variable b1768 : boolean := false;
    variable b1767 : boolean := false;
    variable b1766 : boolean := false;
    variable b1765 : boolean := false;
    variable b1764 : boolean := false;
    variable b1763 : boolean := false;
    variable b1762 : boolean := false;
    variable b1761 : boolean := false;
    variable b1760 : boolean := false;
    variable b1759 : boolean := false;
    variable b1758 : boolean := false;
    variable b1757 : boolean := false;
    variable b1756 : boolean := false;
    variable b1755 : boolean := false;
    variable b1754 : boolean := false;
    variable b1753 : boolean := false;
    variable b1752 : boolean := false;
    variable b1751 : boolean := false;
    variable b1750 : boolean := false;
    variable b1749 : boolean := false;
    variable b1748 : boolean := false;
    variable b1747 : boolean := false;
    variable b1746 : boolean := false;
    variable b1745 : boolean := false;
    variable b1744 : boolean := false;
    variable b1743 : boolean := false;
    variable b1742 : boolean := false;
    variable b1741 : boolean := false;
    variable b1740 : boolean := false;
    variable b1739 : boolean := false;
    variable b1738 : boolean := false;
    variable b1737 : boolean := false;
    variable b1736 : boolean := false;
    variable r1735 : std_logic_vector(0 to 0) := (others => '0');
    variable r1734 : std_logic_vector(0 to 0) := (others => '0');
    variable r1733 : std_logic_vector(0 to 0) := (others => '0');
    variable r1732 : std_logic_vector(0 to 0) := (others => '0');
    variable r1731 : std_logic_vector(0 to 0) := (others => '0');
    variable r1730 : std_logic_vector(0 to 0) := (others => '0');
    variable r1729 : std_logic_vector(0 to 0) := (others => '0');
    variable r1728 : std_logic_vector(0 to 0) := (others => '0');
    variable r1727 : std_logic_vector(0 to 0) := (others => '0');
    variable r1726 : std_logic_vector(0 to 0) := (others => '0');
    variable r1725 : std_logic_vector(0 to 0) := (others => '0');
    variable r1724 : std_logic_vector(0 to 0) := (others => '0');
    variable r1723 : std_logic_vector(0 to 0) := (others => '0');
    variable r1722 : std_logic_vector(0 to 0) := (others => '0');
    variable r1721 : std_logic_vector(0 to 0) := (others => '0');
    variable r1720 : std_logic_vector(0 to 0) := (others => '0');
    variable r1719 : std_logic_vector(0 to 0) := (others => '0');
    variable r1718 : std_logic_vector(0 to 0) := (others => '0');
    variable r1717 : std_logic_vector(0 to 0) := (others => '0');
    variable r1716 : std_logic_vector(0 to 0) := (others => '0');
    variable r1715 : std_logic_vector(0 to 0) := (others => '0');
    variable r1714 : std_logic_vector(0 to 0) := (others => '0');
    variable r1713 : std_logic_vector(0 to 0) := (others => '0');
    variable r1712 : std_logic_vector(0 to 0) := (others => '0');
    variable r1711 : std_logic_vector(0 to 0) := (others => '0');
    variable r1710 : std_logic_vector(0 to 0) := (others => '0');
    variable r1709 : std_logic_vector(0 to 0) := (others => '0');
    variable r1708 : std_logic_vector(0 to 0) := (others => '0');
    variable r1707 : std_logic_vector(0 to 0) := (others => '0');
    variable r1706 : std_logic_vector(0 to 0) := (others => '0');
    variable r1705 : std_logic_vector(0 to 0) := (others => '0');
    variable r1704 : std_logic_vector(0 to 0) := (others => '0');
    variable b1703 : boolean := false;
    variable r1702 : std_logic_vector(0 to 31) := (others => '0');
  begin
    b1703 := true;
    r1704 := r1700(0 to 0);
    r1705 := r1700(1 to 1);
    r1706 := r1700(2 to 2);
    r1707 := r1700(3 to 3);
    r1708 := r1700(4 to 4);
    r1709 := r1700(5 to 5);
    r1710 := r1700(6 to 6);
    r1711 := r1700(7 to 7);
    r1712 := r1700(8 to 8);
    r1713 := r1700(9 to 9);
    r1714 := r1700(10 to 10);
    r1715 := r1700(11 to 11);
    r1716 := r1700(12 to 12);
    r1717 := r1700(13 to 13);
    r1718 := r1700(14 to 14);
    r1719 := r1700(15 to 15);
    r1720 := r1700(16 to 16);
    r1721 := r1700(17 to 17);
    r1722 := r1700(18 to 18);
    r1723 := r1700(19 to 19);
    r1724 := r1700(20 to 20);
    r1725 := r1700(21 to 21);
    r1726 := r1700(22 to 22);
    r1727 := r1700(23 to 23);
    r1728 := r1700(24 to 24);
    r1729 := r1700(25 to 25);
    r1730 := r1700(26 to 26);
    r1731 := r1700(27 to 27);
    r1732 := r1700(28 to 28);
    r1733 := r1700(29 to 29);
    r1734 := r1700(30 to 30);
    r1735 := r1700(31 to 31);
    b1736 := true;
    b1737 := true;
    b1738 := true;
    b1739 := true;
    b1740 := true;
    b1741 := true;
    b1742 := true;
    b1743 := true;
    b1744 := true;
    b1745 := true;
    b1746 := true;
    b1747 := true;
    b1748 := true;
    b1749 := true;
    b1750 := true;
    b1751 := true;
    b1752 := true;
    b1753 := true;
    b1754 := true;
    b1755 := true;
    b1756 := true;
    b1757 := true;
    b1758 := true;
    b1759 := true;
    b1760 := true;
    b1761 := true;
    b1762 := true;
    b1763 := true;
    b1764 := true;
    b1765 := true;
    b1766 := true;
    b1767 := true;
    b1768 := (b1736 AND (b1737 AND (b1738 AND (b1739 AND (b1740 AND (b1741 AND (b1742 AND (b1743 AND (b1744 AND (b1745 AND (b1746 AND (b1747 AND (b1748 AND (b1749 AND (b1750 AND (b1751 AND (b1752 AND (b1753 AND (b1754 AND (b1755 AND (b1756 AND (b1757 AND (b1758 AND (b1759 AND (b1760 AND (b1761 AND (b1762 AND (b1763 AND (b1764 AND (b1765 AND (b1766 AND b1767)))))))))))))))))))))))))))))));
    if b1768 then
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      r1771 := (r1728 & r1729 & r1730 & r1731 & r1732 & r1733 & r1734 & r1735);
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      r1773 := (r1720 & r1721 & r1722 & r1723 & r1724 & r1725 & r1726 & r1727);
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      r1775 := (r1712 & r1713 & r1714 & r1715 & r1716 & r1717 & r1718 & r1719);
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      r1777 := (r1704 & r1705 & r1706 & r1707 & r1708 & r1709 & r1710 & r1711);
      r1778 := (r1771 & r1773 & r1775 & r1777);
      r1702 := r1778;
    end if;
    return r1702;
  end rewire_littleendianp_1699;
  function rewire_sigma3_1533 return std_logic_vector
  is
    variable r1608 : std_logic_vector(0 to 31) := (others => '0');
    variable r1607 : std_logic_vector(0 to 7) := (others => '0');
    variable r1605 : std_logic_vector(0 to 0) := (others => '0');
    variable r1603 : std_logic_vector(0 to 0) := (others => '0');
    variable r1601 : std_logic_vector(0 to 0) := (others => '0');
    variable r1599 : std_logic_vector(0 to 0) := (others => '0');
    variable r1597 : std_logic_vector(0 to 0) := (others => '0');
    variable r1595 : std_logic_vector(0 to 0) := (others => '0');
    variable r1593 : std_logic_vector(0 to 0) := (others => '0');
    variable r1591 : std_logic_vector(0 to 0) := (others => '0');
    variable r1589 : std_logic_vector(0 to 7) := (others => '0');
    variable r1587 : std_logic_vector(0 to 0) := (others => '0');
    variable r1585 : std_logic_vector(0 to 0) := (others => '0');
    variable r1583 : std_logic_vector(0 to 0) := (others => '0');
    variable r1581 : std_logic_vector(0 to 0) := (others => '0');
    variable r1579 : std_logic_vector(0 to 0) := (others => '0');
    variable r1577 : std_logic_vector(0 to 0) := (others => '0');
    variable r1575 : std_logic_vector(0 to 0) := (others => '0');
    variable r1573 : std_logic_vector(0 to 0) := (others => '0');
    variable r1571 : std_logic_vector(0 to 7) := (others => '0');
    variable r1569 : std_logic_vector(0 to 0) := (others => '0');
    variable r1567 : std_logic_vector(0 to 0) := (others => '0');
    variable r1565 : std_logic_vector(0 to 0) := (others => '0');
    variable r1563 : std_logic_vector(0 to 0) := (others => '0');
    variable r1561 : std_logic_vector(0 to 0) := (others => '0');
    variable r1559 : std_logic_vector(0 to 0) := (others => '0');
    variable r1557 : std_logic_vector(0 to 0) := (others => '0');
    variable r1555 : std_logic_vector(0 to 0) := (others => '0');
    variable r1553 : std_logic_vector(0 to 7) := (others => '0');
    variable r1551 : std_logic_vector(0 to 0) := (others => '0');
    variable r1549 : std_logic_vector(0 to 0) := (others => '0');
    variable r1547 : std_logic_vector(0 to 0) := (others => '0');
    variable r1545 : std_logic_vector(0 to 0) := (others => '0');
    variable r1543 : std_logic_vector(0 to 0) := (others => '0');
    variable r1541 : std_logic_vector(0 to 0) := (others => '0');
    variable r1539 : std_logic_vector(0 to 0) := (others => '0');
    variable r1537 : std_logic_vector(0 to 0) := (others => '0');
  begin
    r1537 := "1";
    r1539 := "1";
    r1541 := "0";
    r1543 := "1";
    r1545 := "0";
    r1547 := "0";
    r1549 := "0";
    r1551 := "1";
    r1553 := (r1537 & r1539 & r1541 & r1543 & r1545 & r1547 & r1549 & r1551);
    r1555 := "0";
    r1557 := "1";
    r1559 := "0";
    r1561 := "1";
    r1563 := "1";
    r1565 := "0";
    r1567 := "0";
    r1569 := "1";
    r1571 := (r1555 & r1557 & r1559 & r1561 & r1563 & r1565 & r1567 & r1569);
    r1573 := "1";
    r1575 := "1";
    r1577 := "1";
    r1579 := "1";
    r1581 := "1";
    r1583 := "0";
    r1585 := "1";
    r1587 := "1";
    r1589 := (r1573 & r1575 & r1577 & r1579 & r1581 & r1583 & r1585 & r1587);
    r1591 := "0";
    r1593 := "0";
    r1595 := "1";
    r1597 := "0";
    r1599 := "1";
    r1601 := "0";
    r1603 := "0";
    r1605 := "1";
    r1607 := (r1591 & r1593 & r1595 & r1597 & r1599 & r1601 & r1603 & r1605);
    r1608 := (r1553 & r1571 & r1589 & r1607);
    return r1608;
  end rewire_sigma3_1533;
  function rewire_sigma2_1456 return std_logic_vector
  is
    variable r1531 : std_logic_vector(0 to 31) := (others => '0');
    variable r1530 : std_logic_vector(0 to 7) := (others => '0');
    variable r1528 : std_logic_vector(0 to 0) := (others => '0');
    variable r1526 : std_logic_vector(0 to 0) := (others => '0');
    variable r1524 : std_logic_vector(0 to 0) := (others => '0');
    variable r1522 : std_logic_vector(0 to 0) := (others => '0');
    variable r1520 : std_logic_vector(0 to 0) := (others => '0');
    variable r1518 : std_logic_vector(0 to 0) := (others => '0');
    variable r1516 : std_logic_vector(0 to 0) := (others => '0');
    variable r1514 : std_logic_vector(0 to 0) := (others => '0');
    variable r1512 : std_logic_vector(0 to 7) := (others => '0');
    variable r1510 : std_logic_vector(0 to 0) := (others => '0');
    variable r1508 : std_logic_vector(0 to 0) := (others => '0');
    variable r1506 : std_logic_vector(0 to 0) := (others => '0');
    variable r1504 : std_logic_vector(0 to 0) := (others => '0');
    variable r1502 : std_logic_vector(0 to 0) := (others => '0');
    variable r1500 : std_logic_vector(0 to 0) := (others => '0');
    variable r1498 : std_logic_vector(0 to 0) := (others => '0');
    variable r1496 : std_logic_vector(0 to 0) := (others => '0');
    variable r1494 : std_logic_vector(0 to 7) := (others => '0');
    variable r1492 : std_logic_vector(0 to 0) := (others => '0');
    variable r1490 : std_logic_vector(0 to 0) := (others => '0');
    variable r1488 : std_logic_vector(0 to 0) := (others => '0');
    variable r1486 : std_logic_vector(0 to 0) := (others => '0');
    variable r1484 : std_logic_vector(0 to 0) := (others => '0');
    variable r1482 : std_logic_vector(0 to 0) := (others => '0');
    variable r1480 : std_logic_vector(0 to 0) := (others => '0');
    variable r1478 : std_logic_vector(0 to 0) := (others => '0');
    variable r1476 : std_logic_vector(0 to 7) := (others => '0');
    variable r1474 : std_logic_vector(0 to 0) := (others => '0');
    variable r1472 : std_logic_vector(0 to 0) := (others => '0');
    variable r1470 : std_logic_vector(0 to 0) := (others => '0');
    variable r1468 : std_logic_vector(0 to 0) := (others => '0');
    variable r1466 : std_logic_vector(0 to 0) := (others => '0');
    variable r1464 : std_logic_vector(0 to 0) := (others => '0');
    variable r1462 : std_logic_vector(0 to 0) := (others => '0');
    variable r1460 : std_logic_vector(0 to 0) := (others => '0');
  begin
    r1460 := "1";
    r1462 := "0";
    r1464 := "1";
    r1466 := "1";
    r1468 := "0";
    r1470 := "0";
    r1472 := "1";
    r1474 := "1";
    r1476 := (r1460 & r1462 & r1464 & r1466 & r1468 & r1470 & r1472 & r1474);
    r1478 := "0";
    r1480 := "1";
    r1482 := "0";
    r1484 := "0";
    r1486 := "1";
    r1488 := "0";
    r1490 := "1";
    r1492 := "1";
    r1494 := (r1478 & r1480 & r1482 & r1484 & r1486 & r1488 & r1490 & r1492);
    r1496 := "1";
    r1498 := "0";
    r1500 := "1";
    r1502 := "1";
    r1504 := "1";
    r1506 := "0";
    r1508 := "0";
    r1510 := "1";
    r1512 := (r1496 & r1498 & r1500 & r1502 & r1504 & r1506 & r1508 & r1510);
    r1514 := "0";
    r1516 := "1";
    r1518 := "1";
    r1520 := "0";
    r1522 := "0";
    r1524 := "0";
    r1526 := "0";
    r1528 := "1";
    r1530 := (r1514 & r1516 & r1518 & r1520 & r1522 & r1524 & r1526 & r1528);
    r1531 := (r1476 & r1494 & r1512 & r1530);
    return r1531;
  end rewire_sigma2_1456;
  function rewire_sigma1_1379 return std_logic_vector
  is
    variable r1454 : std_logic_vector(0 to 31) := (others => '0');
    variable r1453 : std_logic_vector(0 to 7) := (others => '0');
    variable r1451 : std_logic_vector(0 to 0) := (others => '0');
    variable r1449 : std_logic_vector(0 to 0) := (others => '0');
    variable r1447 : std_logic_vector(0 to 0) := (others => '0');
    variable r1445 : std_logic_vector(0 to 0) := (others => '0');
    variable r1443 : std_logic_vector(0 to 0) := (others => '0');
    variable r1441 : std_logic_vector(0 to 0) := (others => '0');
    variable r1439 : std_logic_vector(0 to 0) := (others => '0');
    variable r1437 : std_logic_vector(0 to 0) := (others => '0');
    variable r1435 : std_logic_vector(0 to 7) := (others => '0');
    variable r1433 : std_logic_vector(0 to 0) := (others => '0');
    variable r1431 : std_logic_vector(0 to 0) := (others => '0');
    variable r1429 : std_logic_vector(0 to 0) := (others => '0');
    variable r1427 : std_logic_vector(0 to 0) := (others => '0');
    variable r1425 : std_logic_vector(0 to 0) := (others => '0');
    variable r1423 : std_logic_vector(0 to 0) := (others => '0');
    variable r1421 : std_logic_vector(0 to 0) := (others => '0');
    variable r1419 : std_logic_vector(0 to 0) := (others => '0');
    variable r1417 : std_logic_vector(0 to 7) := (others => '0');
    variable r1415 : std_logic_vector(0 to 0) := (others => '0');
    variable r1413 : std_logic_vector(0 to 0) := (others => '0');
    variable r1411 : std_logic_vector(0 to 0) := (others => '0');
    variable r1409 : std_logic_vector(0 to 0) := (others => '0');
    variable r1407 : std_logic_vector(0 to 0) := (others => '0');
    variable r1405 : std_logic_vector(0 to 0) := (others => '0');
    variable r1403 : std_logic_vector(0 to 0) := (others => '0');
    variable r1401 : std_logic_vector(0 to 0) := (others => '0');
    variable r1399 : std_logic_vector(0 to 7) := (others => '0');
    variable r1397 : std_logic_vector(0 to 0) := (others => '0');
    variable r1395 : std_logic_vector(0 to 0) := (others => '0');
    variable r1393 : std_logic_vector(0 to 0) := (others => '0');
    variable r1391 : std_logic_vector(0 to 0) := (others => '0');
    variable r1389 : std_logic_vector(0 to 0) := (others => '0');
    variable r1387 : std_logic_vector(0 to 0) := (others => '0');
    variable r1385 : std_logic_vector(0 to 0) := (others => '0');
    variable r1383 : std_logic_vector(0 to 0) := (others => '0');
  begin
    r1383 := "1";
    r1385 := "0";
    r1387 := "0";
    r1389 := "0";
    r1391 := "1";
    r1393 := "0";
    r1395 := "0";
    r1397 := "1";
    r1399 := (r1383 & r1385 & r1387 & r1389 & r1391 & r1393 & r1395 & r1397);
    r1401 := "1";
    r1403 := "1";
    r1405 := "0";
    r1407 := "1";
    r1409 := "1";
    r1411 := "0";
    r1413 := "0";
    r1415 := "1";
    r1417 := (r1401 & r1403 & r1405 & r1407 & r1409 & r1411 & r1413 & r1415);
    r1419 := "1";
    r1421 := "1";
    r1423 := "1";
    r1425 := "1";
    r1427 := "1";
    r1429 := "0";
    r1431 := "1";
    r1433 := "1";
    r1435 := (r1419 & r1421 & r1423 & r1425 & r1427 & r1429 & r1431 & r1433);
    r1437 := "0";
    r1439 := "0";
    r1441 := "1";
    r1443 := "1";
    r1445 := "0";
    r1447 := "0";
    r1449 := "1";
    r1451 := "1";
    r1453 := (r1437 & r1439 & r1441 & r1443 & r1445 & r1447 & r1449 & r1451);
    r1454 := (r1399 & r1417 & r1435 & r1453);
    return r1454;
  end rewire_sigma1_1379;
  function rewire_sigma0_1302 return std_logic_vector
  is
    variable r1377 : std_logic_vector(0 to 31) := (others => '0');
    variable r1376 : std_logic_vector(0 to 7) := (others => '0');
    variable r1374 : std_logic_vector(0 to 0) := (others => '0');
    variable r1372 : std_logic_vector(0 to 0) := (others => '0');
    variable r1370 : std_logic_vector(0 to 0) := (others => '0');
    variable r1368 : std_logic_vector(0 to 0) := (others => '0');
    variable r1366 : std_logic_vector(0 to 0) := (others => '0');
    variable r1364 : std_logic_vector(0 to 0) := (others => '0');
    variable r1362 : std_logic_vector(0 to 0) := (others => '0');
    variable r1360 : std_logic_vector(0 to 0) := (others => '0');
    variable r1358 : std_logic_vector(0 to 7) := (others => '0');
    variable r1356 : std_logic_vector(0 to 0) := (others => '0');
    variable r1354 : std_logic_vector(0 to 0) := (others => '0');
    variable r1352 : std_logic_vector(0 to 0) := (others => '0');
    variable r1350 : std_logic_vector(0 to 0) := (others => '0');
    variable r1348 : std_logic_vector(0 to 0) := (others => '0');
    variable r1346 : std_logic_vector(0 to 0) := (others => '0');
    variable r1344 : std_logic_vector(0 to 0) := (others => '0');
    variable r1342 : std_logic_vector(0 to 0) := (others => '0');
    variable r1340 : std_logic_vector(0 to 7) := (others => '0');
    variable r1338 : std_logic_vector(0 to 0) := (others => '0');
    variable r1336 : std_logic_vector(0 to 0) := (others => '0');
    variable r1334 : std_logic_vector(0 to 0) := (others => '0');
    variable r1332 : std_logic_vector(0 to 0) := (others => '0');
    variable r1330 : std_logic_vector(0 to 0) := (others => '0');
    variable r1328 : std_logic_vector(0 to 0) := (others => '0');
    variable r1326 : std_logic_vector(0 to 0) := (others => '0');
    variable r1324 : std_logic_vector(0 to 0) := (others => '0');
    variable r1322 : std_logic_vector(0 to 7) := (others => '0');
    variable r1320 : std_logic_vector(0 to 0) := (others => '0');
    variable r1318 : std_logic_vector(0 to 0) := (others => '0');
    variable r1316 : std_logic_vector(0 to 0) := (others => '0');
    variable r1314 : std_logic_vector(0 to 0) := (others => '0');
    variable r1312 : std_logic_vector(0 to 0) := (others => '0');
    variable r1310 : std_logic_vector(0 to 0) := (others => '0');
    variable r1308 : std_logic_vector(0 to 0) := (others => '0');
    variable r1306 : std_logic_vector(0 to 0) := (others => '0');
  begin
    r1306 := "0";
    r1308 := "1";
    r1310 := "0";
    r1312 := "1";
    r1314 := "1";
    r1316 := "0";
    r1318 := "0";
    r1320 := "1";
    r1322 := (r1306 & r1308 & r1310 & r1312 & r1314 & r1316 & r1318 & r1320);
    r1324 := "1";
    r1326 := "1";
    r1328 := "1";
    r1330 := "0";
    r1332 := "0";
    r1334 := "0";
    r1336 := "0";
    r1338 := "1";
    r1340 := (r1324 & r1326 & r1328 & r1330 & r1332 & r1334 & r1336 & r1338);
    r1342 := "1";
    r1344 := "1";
    r1346 := "1";
    r1348 := "1";
    r1350 := "0";
    r1352 := "0";
    r1354 := "0";
    r1356 := "1";
    r1358 := (r1342 & r1344 & r1346 & r1348 & r1350 & r1352 & r1354 & r1356);
    r1360 := "0";
    r1362 := "1";
    r1364 := "1";
    r1366 := "1";
    r1368 := "1";
    r1370 := "0";
    r1372 := "0";
    r1374 := "1";
    r1376 := (r1360 & r1362 & r1364 & r1366 & r1368 & r1370 & r1372 & r1374);
    r1377 := (r1322 & r1340 & r1358 & r1376);
    return r1377;
  end rewire_sigma0_1302;
  function rewire_zerothoutput_3 return std_logic_vector
  is
    variable r1158 : std_logic_vector(0 to 511) := (others => '0');
    variable r1157 : std_logic_vector(0 to 7) := (others => '0');
    variable r1155 : std_logic_vector(0 to 0) := (others => '0');
    variable r1153 : std_logic_vector(0 to 0) := (others => '0');
    variable r1151 : std_logic_vector(0 to 0) := (others => '0');
    variable r1149 : std_logic_vector(0 to 0) := (others => '0');
    variable r1147 : std_logic_vector(0 to 0) := (others => '0');
    variable r1145 : std_logic_vector(0 to 0) := (others => '0');
    variable r1143 : std_logic_vector(0 to 0) := (others => '0');
    variable r1141 : std_logic_vector(0 to 0) := (others => '0');
    variable r1139 : std_logic_vector(0 to 7) := (others => '0');
    variable r1137 : std_logic_vector(0 to 0) := (others => '0');
    variable r1135 : std_logic_vector(0 to 0) := (others => '0');
    variable r1133 : std_logic_vector(0 to 0) := (others => '0');
    variable r1131 : std_logic_vector(0 to 0) := (others => '0');
    variable r1129 : std_logic_vector(0 to 0) := (others => '0');
    variable r1127 : std_logic_vector(0 to 0) := (others => '0');
    variable r1125 : std_logic_vector(0 to 0) := (others => '0');
    variable r1123 : std_logic_vector(0 to 0) := (others => '0');
    variable r1121 : std_logic_vector(0 to 7) := (others => '0');
    variable r1119 : std_logic_vector(0 to 0) := (others => '0');
    variable r1117 : std_logic_vector(0 to 0) := (others => '0');
    variable r1115 : std_logic_vector(0 to 0) := (others => '0');
    variable r1113 : std_logic_vector(0 to 0) := (others => '0');
    variable r1111 : std_logic_vector(0 to 0) := (others => '0');
    variable r1109 : std_logic_vector(0 to 0) := (others => '0');
    variable r1107 : std_logic_vector(0 to 0) := (others => '0');
    variable r1105 : std_logic_vector(0 to 0) := (others => '0');
    variable r1103 : std_logic_vector(0 to 7) := (others => '0');
    variable r1101 : std_logic_vector(0 to 0) := (others => '0');
    variable r1099 : std_logic_vector(0 to 0) := (others => '0');
    variable r1097 : std_logic_vector(0 to 0) := (others => '0');
    variable r1095 : std_logic_vector(0 to 0) := (others => '0');
    variable r1093 : std_logic_vector(0 to 0) := (others => '0');
    variable r1091 : std_logic_vector(0 to 0) := (others => '0');
    variable r1089 : std_logic_vector(0 to 0) := (others => '0');
    variable r1087 : std_logic_vector(0 to 0) := (others => '0');
    variable r1085 : std_logic_vector(0 to 7) := (others => '0');
    variable r1083 : std_logic_vector(0 to 0) := (others => '0');
    variable r1081 : std_logic_vector(0 to 0) := (others => '0');
    variable r1079 : std_logic_vector(0 to 0) := (others => '0');
    variable r1077 : std_logic_vector(0 to 0) := (others => '0');
    variable r1075 : std_logic_vector(0 to 0) := (others => '0');
    variable r1073 : std_logic_vector(0 to 0) := (others => '0');
    variable r1071 : std_logic_vector(0 to 0) := (others => '0');
    variable r1069 : std_logic_vector(0 to 0) := (others => '0');
    variable r1067 : std_logic_vector(0 to 7) := (others => '0');
    variable r1065 : std_logic_vector(0 to 0) := (others => '0');
    variable r1063 : std_logic_vector(0 to 0) := (others => '0');
    variable r1061 : std_logic_vector(0 to 0) := (others => '0');
    variable r1059 : std_logic_vector(0 to 0) := (others => '0');
    variable r1057 : std_logic_vector(0 to 0) := (others => '0');
    variable r1055 : std_logic_vector(0 to 0) := (others => '0');
    variable r1053 : std_logic_vector(0 to 0) := (others => '0');
    variable r1051 : std_logic_vector(0 to 0) := (others => '0');
    variable r1049 : std_logic_vector(0 to 7) := (others => '0');
    variable r1047 : std_logic_vector(0 to 0) := (others => '0');
    variable r1045 : std_logic_vector(0 to 0) := (others => '0');
    variable r1043 : std_logic_vector(0 to 0) := (others => '0');
    variable r1041 : std_logic_vector(0 to 0) := (others => '0');
    variable r1039 : std_logic_vector(0 to 0) := (others => '0');
    variable r1037 : std_logic_vector(0 to 0) := (others => '0');
    variable r1035 : std_logic_vector(0 to 0) := (others => '0');
    variable r1033 : std_logic_vector(0 to 0) := (others => '0');
    variable r1031 : std_logic_vector(0 to 7) := (others => '0');
    variable r1029 : std_logic_vector(0 to 0) := (others => '0');
    variable r1027 : std_logic_vector(0 to 0) := (others => '0');
    variable r1025 : std_logic_vector(0 to 0) := (others => '0');
    variable r1023 : std_logic_vector(0 to 0) := (others => '0');
    variable r1021 : std_logic_vector(0 to 0) := (others => '0');
    variable r1019 : std_logic_vector(0 to 0) := (others => '0');
    variable r1017 : std_logic_vector(0 to 0) := (others => '0');
    variable r1015 : std_logic_vector(0 to 0) := (others => '0');
    variable r1013 : std_logic_vector(0 to 7) := (others => '0');
    variable r1011 : std_logic_vector(0 to 0) := (others => '0');
    variable r1009 : std_logic_vector(0 to 0) := (others => '0');
    variable r1007 : std_logic_vector(0 to 0) := (others => '0');
    variable r1005 : std_logic_vector(0 to 0) := (others => '0');
    variable r1003 : std_logic_vector(0 to 0) := (others => '0');
    variable r1001 : std_logic_vector(0 to 0) := (others => '0');
    variable r999 : std_logic_vector(0 to 0) := (others => '0');
    variable r997 : std_logic_vector(0 to 0) := (others => '0');
    variable r995 : std_logic_vector(0 to 7) := (others => '0');
    variable r993 : std_logic_vector(0 to 0) := (others => '0');
    variable r991 : std_logic_vector(0 to 0) := (others => '0');
    variable r989 : std_logic_vector(0 to 0) := (others => '0');
    variable r987 : std_logic_vector(0 to 0) := (others => '0');
    variable r985 : std_logic_vector(0 to 0) := (others => '0');
    variable r983 : std_logic_vector(0 to 0) := (others => '0');
    variable r981 : std_logic_vector(0 to 0) := (others => '0');
    variable r979 : std_logic_vector(0 to 0) := (others => '0');
    variable r977 : std_logic_vector(0 to 7) := (others => '0');
    variable r975 : std_logic_vector(0 to 0) := (others => '0');
    variable r973 : std_logic_vector(0 to 0) := (others => '0');
    variable r971 : std_logic_vector(0 to 0) := (others => '0');
    variable r969 : std_logic_vector(0 to 0) := (others => '0');
    variable r967 : std_logic_vector(0 to 0) := (others => '0');
    variable r965 : std_logic_vector(0 to 0) := (others => '0');
    variable r963 : std_logic_vector(0 to 0) := (others => '0');
    variable r961 : std_logic_vector(0 to 0) := (others => '0');
    variable r959 : std_logic_vector(0 to 7) := (others => '0');
    variable r957 : std_logic_vector(0 to 0) := (others => '0');
    variable r955 : std_logic_vector(0 to 0) := (others => '0');
    variable r953 : std_logic_vector(0 to 0) := (others => '0');
    variable r951 : std_logic_vector(0 to 0) := (others => '0');
    variable r949 : std_logic_vector(0 to 0) := (others => '0');
    variable r947 : std_logic_vector(0 to 0) := (others => '0');
    variable r945 : std_logic_vector(0 to 0) := (others => '0');
    variable r943 : std_logic_vector(0 to 0) := (others => '0');
    variable r941 : std_logic_vector(0 to 7) := (others => '0');
    variable r939 : std_logic_vector(0 to 0) := (others => '0');
    variable r937 : std_logic_vector(0 to 0) := (others => '0');
    variable r935 : std_logic_vector(0 to 0) := (others => '0');
    variable r933 : std_logic_vector(0 to 0) := (others => '0');
    variable r931 : std_logic_vector(0 to 0) := (others => '0');
    variable r929 : std_logic_vector(0 to 0) := (others => '0');
    variable r927 : std_logic_vector(0 to 0) := (others => '0');
    variable r925 : std_logic_vector(0 to 0) := (others => '0');
    variable r923 : std_logic_vector(0 to 7) := (others => '0');
    variable r921 : std_logic_vector(0 to 0) := (others => '0');
    variable r919 : std_logic_vector(0 to 0) := (others => '0');
    variable r917 : std_logic_vector(0 to 0) := (others => '0');
    variable r915 : std_logic_vector(0 to 0) := (others => '0');
    variable r913 : std_logic_vector(0 to 0) := (others => '0');
    variable r911 : std_logic_vector(0 to 0) := (others => '0');
    variable r909 : std_logic_vector(0 to 0) := (others => '0');
    variable r907 : std_logic_vector(0 to 0) := (others => '0');
    variable r905 : std_logic_vector(0 to 7) := (others => '0');
    variable r903 : std_logic_vector(0 to 0) := (others => '0');
    variable r901 : std_logic_vector(0 to 0) := (others => '0');
    variable r899 : std_logic_vector(0 to 0) := (others => '0');
    variable r897 : std_logic_vector(0 to 0) := (others => '0');
    variable r895 : std_logic_vector(0 to 0) := (others => '0');
    variable r893 : std_logic_vector(0 to 0) := (others => '0');
    variable r891 : std_logic_vector(0 to 0) := (others => '0');
    variable r889 : std_logic_vector(0 to 0) := (others => '0');
    variable r887 : std_logic_vector(0 to 7) := (others => '0');
    variable r885 : std_logic_vector(0 to 0) := (others => '0');
    variable r883 : std_logic_vector(0 to 0) := (others => '0');
    variable r881 : std_logic_vector(0 to 0) := (others => '0');
    variable r879 : std_logic_vector(0 to 0) := (others => '0');
    variable r877 : std_logic_vector(0 to 0) := (others => '0');
    variable r875 : std_logic_vector(0 to 0) := (others => '0');
    variable r873 : std_logic_vector(0 to 0) := (others => '0');
    variable r871 : std_logic_vector(0 to 0) := (others => '0');
    variable r869 : std_logic_vector(0 to 7) := (others => '0');
    variable r867 : std_logic_vector(0 to 0) := (others => '0');
    variable r865 : std_logic_vector(0 to 0) := (others => '0');
    variable r863 : std_logic_vector(0 to 0) := (others => '0');
    variable r861 : std_logic_vector(0 to 0) := (others => '0');
    variable r859 : std_logic_vector(0 to 0) := (others => '0');
    variable r857 : std_logic_vector(0 to 0) := (others => '0');
    variable r855 : std_logic_vector(0 to 0) := (others => '0');
    variable r853 : std_logic_vector(0 to 0) := (others => '0');
    variable r851 : std_logic_vector(0 to 7) := (others => '0');
    variable r849 : std_logic_vector(0 to 0) := (others => '0');
    variable r847 : std_logic_vector(0 to 0) := (others => '0');
    variable r845 : std_logic_vector(0 to 0) := (others => '0');
    variable r843 : std_logic_vector(0 to 0) := (others => '0');
    variable r841 : std_logic_vector(0 to 0) := (others => '0');
    variable r839 : std_logic_vector(0 to 0) := (others => '0');
    variable r837 : std_logic_vector(0 to 0) := (others => '0');
    variable r835 : std_logic_vector(0 to 0) := (others => '0');
    variable r833 : std_logic_vector(0 to 7) := (others => '0');
    variable r831 : std_logic_vector(0 to 0) := (others => '0');
    variable r829 : std_logic_vector(0 to 0) := (others => '0');
    variable r827 : std_logic_vector(0 to 0) := (others => '0');
    variable r825 : std_logic_vector(0 to 0) := (others => '0');
    variable r823 : std_logic_vector(0 to 0) := (others => '0');
    variable r821 : std_logic_vector(0 to 0) := (others => '0');
    variable r819 : std_logic_vector(0 to 0) := (others => '0');
    variable r817 : std_logic_vector(0 to 0) := (others => '0');
    variable r815 : std_logic_vector(0 to 7) := (others => '0');
    variable r813 : std_logic_vector(0 to 0) := (others => '0');
    variable r811 : std_logic_vector(0 to 0) := (others => '0');
    variable r809 : std_logic_vector(0 to 0) := (others => '0');
    variable r807 : std_logic_vector(0 to 0) := (others => '0');
    variable r805 : std_logic_vector(0 to 0) := (others => '0');
    variable r803 : std_logic_vector(0 to 0) := (others => '0');
    variable r801 : std_logic_vector(0 to 0) := (others => '0');
    variable r799 : std_logic_vector(0 to 0) := (others => '0');
    variable r797 : std_logic_vector(0 to 7) := (others => '0');
    variable r795 : std_logic_vector(0 to 0) := (others => '0');
    variable r793 : std_logic_vector(0 to 0) := (others => '0');
    variable r791 : std_logic_vector(0 to 0) := (others => '0');
    variable r789 : std_logic_vector(0 to 0) := (others => '0');
    variable r787 : std_logic_vector(0 to 0) := (others => '0');
    variable r785 : std_logic_vector(0 to 0) := (others => '0');
    variable r783 : std_logic_vector(0 to 0) := (others => '0');
    variable r781 : std_logic_vector(0 to 0) := (others => '0');
    variable r779 : std_logic_vector(0 to 7) := (others => '0');
    variable r777 : std_logic_vector(0 to 0) := (others => '0');
    variable r775 : std_logic_vector(0 to 0) := (others => '0');
    variable r773 : std_logic_vector(0 to 0) := (others => '0');
    variable r771 : std_logic_vector(0 to 0) := (others => '0');
    variable r769 : std_logic_vector(0 to 0) := (others => '0');
    variable r767 : std_logic_vector(0 to 0) := (others => '0');
    variable r765 : std_logic_vector(0 to 0) := (others => '0');
    variable r763 : std_logic_vector(0 to 0) := (others => '0');
    variable r761 : std_logic_vector(0 to 7) := (others => '0');
    variable r759 : std_logic_vector(0 to 0) := (others => '0');
    variable r757 : std_logic_vector(0 to 0) := (others => '0');
    variable r755 : std_logic_vector(0 to 0) := (others => '0');
    variable r753 : std_logic_vector(0 to 0) := (others => '0');
    variable r751 : std_logic_vector(0 to 0) := (others => '0');
    variable r749 : std_logic_vector(0 to 0) := (others => '0');
    variable r747 : std_logic_vector(0 to 0) := (others => '0');
    variable r745 : std_logic_vector(0 to 0) := (others => '0');
    variable r743 : std_logic_vector(0 to 7) := (others => '0');
    variable r741 : std_logic_vector(0 to 0) := (others => '0');
    variable r739 : std_logic_vector(0 to 0) := (others => '0');
    variable r737 : std_logic_vector(0 to 0) := (others => '0');
    variable r735 : std_logic_vector(0 to 0) := (others => '0');
    variable r733 : std_logic_vector(0 to 0) := (others => '0');
    variable r731 : std_logic_vector(0 to 0) := (others => '0');
    variable r729 : std_logic_vector(0 to 0) := (others => '0');
    variable r727 : std_logic_vector(0 to 0) := (others => '0');
    variable r725 : std_logic_vector(0 to 7) := (others => '0');
    variable r723 : std_logic_vector(0 to 0) := (others => '0');
    variable r721 : std_logic_vector(0 to 0) := (others => '0');
    variable r719 : std_logic_vector(0 to 0) := (others => '0');
    variable r717 : std_logic_vector(0 to 0) := (others => '0');
    variable r715 : std_logic_vector(0 to 0) := (others => '0');
    variable r713 : std_logic_vector(0 to 0) := (others => '0');
    variable r711 : std_logic_vector(0 to 0) := (others => '0');
    variable r709 : std_logic_vector(0 to 0) := (others => '0');
    variable r707 : std_logic_vector(0 to 7) := (others => '0');
    variable r705 : std_logic_vector(0 to 0) := (others => '0');
    variable r703 : std_logic_vector(0 to 0) := (others => '0');
    variable r701 : std_logic_vector(0 to 0) := (others => '0');
    variable r699 : std_logic_vector(0 to 0) := (others => '0');
    variable r697 : std_logic_vector(0 to 0) := (others => '0');
    variable r695 : std_logic_vector(0 to 0) := (others => '0');
    variable r693 : std_logic_vector(0 to 0) := (others => '0');
    variable r691 : std_logic_vector(0 to 0) := (others => '0');
    variable r689 : std_logic_vector(0 to 7) := (others => '0');
    variable r687 : std_logic_vector(0 to 0) := (others => '0');
    variable r685 : std_logic_vector(0 to 0) := (others => '0');
    variable r683 : std_logic_vector(0 to 0) := (others => '0');
    variable r681 : std_logic_vector(0 to 0) := (others => '0');
    variable r679 : std_logic_vector(0 to 0) := (others => '0');
    variable r677 : std_logic_vector(0 to 0) := (others => '0');
    variable r675 : std_logic_vector(0 to 0) := (others => '0');
    variable r673 : std_logic_vector(0 to 0) := (others => '0');
    variable r671 : std_logic_vector(0 to 7) := (others => '0');
    variable r669 : std_logic_vector(0 to 0) := (others => '0');
    variable r667 : std_logic_vector(0 to 0) := (others => '0');
    variable r665 : std_logic_vector(0 to 0) := (others => '0');
    variable r663 : std_logic_vector(0 to 0) := (others => '0');
    variable r661 : std_logic_vector(0 to 0) := (others => '0');
    variable r659 : std_logic_vector(0 to 0) := (others => '0');
    variable r657 : std_logic_vector(0 to 0) := (others => '0');
    variable r655 : std_logic_vector(0 to 0) := (others => '0');
    variable r653 : std_logic_vector(0 to 7) := (others => '0');
    variable r651 : std_logic_vector(0 to 0) := (others => '0');
    variable r649 : std_logic_vector(0 to 0) := (others => '0');
    variable r647 : std_logic_vector(0 to 0) := (others => '0');
    variable r645 : std_logic_vector(0 to 0) := (others => '0');
    variable r643 : std_logic_vector(0 to 0) := (others => '0');
    variable r641 : std_logic_vector(0 to 0) := (others => '0');
    variable r639 : std_logic_vector(0 to 0) := (others => '0');
    variable r637 : std_logic_vector(0 to 0) := (others => '0');
    variable r635 : std_logic_vector(0 to 7) := (others => '0');
    variable r633 : std_logic_vector(0 to 0) := (others => '0');
    variable r631 : std_logic_vector(0 to 0) := (others => '0');
    variable r629 : std_logic_vector(0 to 0) := (others => '0');
    variable r627 : std_logic_vector(0 to 0) := (others => '0');
    variable r625 : std_logic_vector(0 to 0) := (others => '0');
    variable r623 : std_logic_vector(0 to 0) := (others => '0');
    variable r621 : std_logic_vector(0 to 0) := (others => '0');
    variable r619 : std_logic_vector(0 to 0) := (others => '0');
    variable r617 : std_logic_vector(0 to 7) := (others => '0');
    variable r615 : std_logic_vector(0 to 0) := (others => '0');
    variable r613 : std_logic_vector(0 to 0) := (others => '0');
    variable r611 : std_logic_vector(0 to 0) := (others => '0');
    variable r609 : std_logic_vector(0 to 0) := (others => '0');
    variable r607 : std_logic_vector(0 to 0) := (others => '0');
    variable r605 : std_logic_vector(0 to 0) := (others => '0');
    variable r603 : std_logic_vector(0 to 0) := (others => '0');
    variable r601 : std_logic_vector(0 to 0) := (others => '0');
    variable r599 : std_logic_vector(0 to 7) := (others => '0');
    variable r597 : std_logic_vector(0 to 0) := (others => '0');
    variable r595 : std_logic_vector(0 to 0) := (others => '0');
    variable r593 : std_logic_vector(0 to 0) := (others => '0');
    variable r591 : std_logic_vector(0 to 0) := (others => '0');
    variable r589 : std_logic_vector(0 to 0) := (others => '0');
    variable r587 : std_logic_vector(0 to 0) := (others => '0');
    variable r585 : std_logic_vector(0 to 0) := (others => '0');
    variable r583 : std_logic_vector(0 to 0) := (others => '0');
    variable r581 : std_logic_vector(0 to 7) := (others => '0');
    variable r579 : std_logic_vector(0 to 0) := (others => '0');
    variable r577 : std_logic_vector(0 to 0) := (others => '0');
    variable r575 : std_logic_vector(0 to 0) := (others => '0');
    variable r573 : std_logic_vector(0 to 0) := (others => '0');
    variable r571 : std_logic_vector(0 to 0) := (others => '0');
    variable r569 : std_logic_vector(0 to 0) := (others => '0');
    variable r567 : std_logic_vector(0 to 0) := (others => '0');
    variable r565 : std_logic_vector(0 to 0) := (others => '0');
    variable r563 : std_logic_vector(0 to 7) := (others => '0');
    variable r561 : std_logic_vector(0 to 0) := (others => '0');
    variable r559 : std_logic_vector(0 to 0) := (others => '0');
    variable r557 : std_logic_vector(0 to 0) := (others => '0');
    variable r555 : std_logic_vector(0 to 0) := (others => '0');
    variable r553 : std_logic_vector(0 to 0) := (others => '0');
    variable r551 : std_logic_vector(0 to 0) := (others => '0');
    variable r549 : std_logic_vector(0 to 0) := (others => '0');
    variable r547 : std_logic_vector(0 to 0) := (others => '0');
    variable r545 : std_logic_vector(0 to 7) := (others => '0');
    variable r543 : std_logic_vector(0 to 0) := (others => '0');
    variable r541 : std_logic_vector(0 to 0) := (others => '0');
    variable r539 : std_logic_vector(0 to 0) := (others => '0');
    variable r537 : std_logic_vector(0 to 0) := (others => '0');
    variable r535 : std_logic_vector(0 to 0) := (others => '0');
    variable r533 : std_logic_vector(0 to 0) := (others => '0');
    variable r531 : std_logic_vector(0 to 0) := (others => '0');
    variable r529 : std_logic_vector(0 to 0) := (others => '0');
    variable r527 : std_logic_vector(0 to 7) := (others => '0');
    variable r525 : std_logic_vector(0 to 0) := (others => '0');
    variable r523 : std_logic_vector(0 to 0) := (others => '0');
    variable r521 : std_logic_vector(0 to 0) := (others => '0');
    variable r519 : std_logic_vector(0 to 0) := (others => '0');
    variable r517 : std_logic_vector(0 to 0) := (others => '0');
    variable r515 : std_logic_vector(0 to 0) := (others => '0');
    variable r513 : std_logic_vector(0 to 0) := (others => '0');
    variable r511 : std_logic_vector(0 to 0) := (others => '0');
    variable r509 : std_logic_vector(0 to 7) := (others => '0');
    variable r507 : std_logic_vector(0 to 0) := (others => '0');
    variable r505 : std_logic_vector(0 to 0) := (others => '0');
    variable r503 : std_logic_vector(0 to 0) := (others => '0');
    variable r501 : std_logic_vector(0 to 0) := (others => '0');
    variable r499 : std_logic_vector(0 to 0) := (others => '0');
    variable r497 : std_logic_vector(0 to 0) := (others => '0');
    variable r495 : std_logic_vector(0 to 0) := (others => '0');
    variable r493 : std_logic_vector(0 to 0) := (others => '0');
    variable r491 : std_logic_vector(0 to 7) := (others => '0');
    variable r489 : std_logic_vector(0 to 0) := (others => '0');
    variable r487 : std_logic_vector(0 to 0) := (others => '0');
    variable r485 : std_logic_vector(0 to 0) := (others => '0');
    variable r483 : std_logic_vector(0 to 0) := (others => '0');
    variable r481 : std_logic_vector(0 to 0) := (others => '0');
    variable r479 : std_logic_vector(0 to 0) := (others => '0');
    variable r477 : std_logic_vector(0 to 0) := (others => '0');
    variable r475 : std_logic_vector(0 to 0) := (others => '0');
    variable r473 : std_logic_vector(0 to 7) := (others => '0');
    variable r471 : std_logic_vector(0 to 0) := (others => '0');
    variable r469 : std_logic_vector(0 to 0) := (others => '0');
    variable r467 : std_logic_vector(0 to 0) := (others => '0');
    variable r465 : std_logic_vector(0 to 0) := (others => '0');
    variable r463 : std_logic_vector(0 to 0) := (others => '0');
    variable r461 : std_logic_vector(0 to 0) := (others => '0');
    variable r459 : std_logic_vector(0 to 0) := (others => '0');
    variable r457 : std_logic_vector(0 to 0) := (others => '0');
    variable r455 : std_logic_vector(0 to 7) := (others => '0');
    variable r453 : std_logic_vector(0 to 0) := (others => '0');
    variable r451 : std_logic_vector(0 to 0) := (others => '0');
    variable r449 : std_logic_vector(0 to 0) := (others => '0');
    variable r447 : std_logic_vector(0 to 0) := (others => '0');
    variable r445 : std_logic_vector(0 to 0) := (others => '0');
    variable r443 : std_logic_vector(0 to 0) := (others => '0');
    variable r441 : std_logic_vector(0 to 0) := (others => '0');
    variable r439 : std_logic_vector(0 to 0) := (others => '0');
    variable r437 : std_logic_vector(0 to 7) := (others => '0');
    variable r435 : std_logic_vector(0 to 0) := (others => '0');
    variable r433 : std_logic_vector(0 to 0) := (others => '0');
    variable r431 : std_logic_vector(0 to 0) := (others => '0');
    variable r429 : std_logic_vector(0 to 0) := (others => '0');
    variable r427 : std_logic_vector(0 to 0) := (others => '0');
    variable r425 : std_logic_vector(0 to 0) := (others => '0');
    variable r423 : std_logic_vector(0 to 0) := (others => '0');
    variable r421 : std_logic_vector(0 to 0) := (others => '0');
    variable r419 : std_logic_vector(0 to 7) := (others => '0');
    variable r417 : std_logic_vector(0 to 0) := (others => '0');
    variable r415 : std_logic_vector(0 to 0) := (others => '0');
    variable r413 : std_logic_vector(0 to 0) := (others => '0');
    variable r411 : std_logic_vector(0 to 0) := (others => '0');
    variable r409 : std_logic_vector(0 to 0) := (others => '0');
    variable r407 : std_logic_vector(0 to 0) := (others => '0');
    variable r405 : std_logic_vector(0 to 0) := (others => '0');
    variable r403 : std_logic_vector(0 to 0) := (others => '0');
    variable r401 : std_logic_vector(0 to 7) := (others => '0');
    variable r399 : std_logic_vector(0 to 0) := (others => '0');
    variable r397 : std_logic_vector(0 to 0) := (others => '0');
    variable r395 : std_logic_vector(0 to 0) := (others => '0');
    variable r393 : std_logic_vector(0 to 0) := (others => '0');
    variable r391 : std_logic_vector(0 to 0) := (others => '0');
    variable r389 : std_logic_vector(0 to 0) := (others => '0');
    variable r387 : std_logic_vector(0 to 0) := (others => '0');
    variable r385 : std_logic_vector(0 to 0) := (others => '0');
    variable r383 : std_logic_vector(0 to 7) := (others => '0');
    variable r381 : std_logic_vector(0 to 0) := (others => '0');
    variable r379 : std_logic_vector(0 to 0) := (others => '0');
    variable r377 : std_logic_vector(0 to 0) := (others => '0');
    variable r375 : std_logic_vector(0 to 0) := (others => '0');
    variable r373 : std_logic_vector(0 to 0) := (others => '0');
    variable r371 : std_logic_vector(0 to 0) := (others => '0');
    variable r369 : std_logic_vector(0 to 0) := (others => '0');
    variable r367 : std_logic_vector(0 to 0) := (others => '0');
    variable r365 : std_logic_vector(0 to 7) := (others => '0');
    variable r363 : std_logic_vector(0 to 0) := (others => '0');
    variable r361 : std_logic_vector(0 to 0) := (others => '0');
    variable r359 : std_logic_vector(0 to 0) := (others => '0');
    variable r357 : std_logic_vector(0 to 0) := (others => '0');
    variable r355 : std_logic_vector(0 to 0) := (others => '0');
    variable r353 : std_logic_vector(0 to 0) := (others => '0');
    variable r351 : std_logic_vector(0 to 0) := (others => '0');
    variable r349 : std_logic_vector(0 to 0) := (others => '0');
    variable r347 : std_logic_vector(0 to 7) := (others => '0');
    variable r345 : std_logic_vector(0 to 0) := (others => '0');
    variable r343 : std_logic_vector(0 to 0) := (others => '0');
    variable r341 : std_logic_vector(0 to 0) := (others => '0');
    variable r339 : std_logic_vector(0 to 0) := (others => '0');
    variable r337 : std_logic_vector(0 to 0) := (others => '0');
    variable r335 : std_logic_vector(0 to 0) := (others => '0');
    variable r333 : std_logic_vector(0 to 0) := (others => '0');
    variable r331 : std_logic_vector(0 to 0) := (others => '0');
    variable r329 : std_logic_vector(0 to 7) := (others => '0');
    variable r327 : std_logic_vector(0 to 0) := (others => '0');
    variable r325 : std_logic_vector(0 to 0) := (others => '0');
    variable r323 : std_logic_vector(0 to 0) := (others => '0');
    variable r321 : std_logic_vector(0 to 0) := (others => '0');
    variable r319 : std_logic_vector(0 to 0) := (others => '0');
    variable r317 : std_logic_vector(0 to 0) := (others => '0');
    variable r315 : std_logic_vector(0 to 0) := (others => '0');
    variable r313 : std_logic_vector(0 to 0) := (others => '0');
    variable r311 : std_logic_vector(0 to 7) := (others => '0');
    variable r309 : std_logic_vector(0 to 0) := (others => '0');
    variable r307 : std_logic_vector(0 to 0) := (others => '0');
    variable r305 : std_logic_vector(0 to 0) := (others => '0');
    variable r303 : std_logic_vector(0 to 0) := (others => '0');
    variable r301 : std_logic_vector(0 to 0) := (others => '0');
    variable r299 : std_logic_vector(0 to 0) := (others => '0');
    variable r297 : std_logic_vector(0 to 0) := (others => '0');
    variable r295 : std_logic_vector(0 to 0) := (others => '0');
    variable r293 : std_logic_vector(0 to 7) := (others => '0');
    variable r291 : std_logic_vector(0 to 0) := (others => '0');
    variable r289 : std_logic_vector(0 to 0) := (others => '0');
    variable r287 : std_logic_vector(0 to 0) := (others => '0');
    variable r285 : std_logic_vector(0 to 0) := (others => '0');
    variable r283 : std_logic_vector(0 to 0) := (others => '0');
    variable r281 : std_logic_vector(0 to 0) := (others => '0');
    variable r279 : std_logic_vector(0 to 0) := (others => '0');
    variable r277 : std_logic_vector(0 to 0) := (others => '0');
    variable r275 : std_logic_vector(0 to 7) := (others => '0');
    variable r273 : std_logic_vector(0 to 0) := (others => '0');
    variable r271 : std_logic_vector(0 to 0) := (others => '0');
    variable r269 : std_logic_vector(0 to 0) := (others => '0');
    variable r267 : std_logic_vector(0 to 0) := (others => '0');
    variable r265 : std_logic_vector(0 to 0) := (others => '0');
    variable r263 : std_logic_vector(0 to 0) := (others => '0');
    variable r261 : std_logic_vector(0 to 0) := (others => '0');
    variable r259 : std_logic_vector(0 to 0) := (others => '0');
    variable r257 : std_logic_vector(0 to 7) := (others => '0');
    variable r255 : std_logic_vector(0 to 0) := (others => '0');
    variable r253 : std_logic_vector(0 to 0) := (others => '0');
    variable r251 : std_logic_vector(0 to 0) := (others => '0');
    variable r249 : std_logic_vector(0 to 0) := (others => '0');
    variable r247 : std_logic_vector(0 to 0) := (others => '0');
    variable r245 : std_logic_vector(0 to 0) := (others => '0');
    variable r243 : std_logic_vector(0 to 0) := (others => '0');
    variable r241 : std_logic_vector(0 to 0) := (others => '0');
    variable r239 : std_logic_vector(0 to 7) := (others => '0');
    variable r237 : std_logic_vector(0 to 0) := (others => '0');
    variable r235 : std_logic_vector(0 to 0) := (others => '0');
    variable r233 : std_logic_vector(0 to 0) := (others => '0');
    variable r231 : std_logic_vector(0 to 0) := (others => '0');
    variable r229 : std_logic_vector(0 to 0) := (others => '0');
    variable r227 : std_logic_vector(0 to 0) := (others => '0');
    variable r225 : std_logic_vector(0 to 0) := (others => '0');
    variable r223 : std_logic_vector(0 to 0) := (others => '0');
    variable r221 : std_logic_vector(0 to 7) := (others => '0');
    variable r219 : std_logic_vector(0 to 0) := (others => '0');
    variable r217 : std_logic_vector(0 to 0) := (others => '0');
    variable r215 : std_logic_vector(0 to 0) := (others => '0');
    variable r213 : std_logic_vector(0 to 0) := (others => '0');
    variable r211 : std_logic_vector(0 to 0) := (others => '0');
    variable r209 : std_logic_vector(0 to 0) := (others => '0');
    variable r207 : std_logic_vector(0 to 0) := (others => '0');
    variable r205 : std_logic_vector(0 to 0) := (others => '0');
    variable r203 : std_logic_vector(0 to 7) := (others => '0');
    variable r201 : std_logic_vector(0 to 0) := (others => '0');
    variable r199 : std_logic_vector(0 to 0) := (others => '0');
    variable r197 : std_logic_vector(0 to 0) := (others => '0');
    variable r195 : std_logic_vector(0 to 0) := (others => '0');
    variable r193 : std_logic_vector(0 to 0) := (others => '0');
    variable r191 : std_logic_vector(0 to 0) := (others => '0');
    variable r189 : std_logic_vector(0 to 0) := (others => '0');
    variable r187 : std_logic_vector(0 to 0) := (others => '0');
    variable r185 : std_logic_vector(0 to 7) := (others => '0');
    variable r183 : std_logic_vector(0 to 0) := (others => '0');
    variable r181 : std_logic_vector(0 to 0) := (others => '0');
    variable r179 : std_logic_vector(0 to 0) := (others => '0');
    variable r177 : std_logic_vector(0 to 0) := (others => '0');
    variable r175 : std_logic_vector(0 to 0) := (others => '0');
    variable r173 : std_logic_vector(0 to 0) := (others => '0');
    variable r171 : std_logic_vector(0 to 0) := (others => '0');
    variable r169 : std_logic_vector(0 to 0) := (others => '0');
    variable r167 : std_logic_vector(0 to 7) := (others => '0');
    variable r165 : std_logic_vector(0 to 0) := (others => '0');
    variable r163 : std_logic_vector(0 to 0) := (others => '0');
    variable r161 : std_logic_vector(0 to 0) := (others => '0');
    variable r159 : std_logic_vector(0 to 0) := (others => '0');
    variable r157 : std_logic_vector(0 to 0) := (others => '0');
    variable r155 : std_logic_vector(0 to 0) := (others => '0');
    variable r153 : std_logic_vector(0 to 0) := (others => '0');
    variable r151 : std_logic_vector(0 to 0) := (others => '0');
    variable r149 : std_logic_vector(0 to 7) := (others => '0');
    variable r147 : std_logic_vector(0 to 0) := (others => '0');
    variable r145 : std_logic_vector(0 to 0) := (others => '0');
    variable r143 : std_logic_vector(0 to 0) := (others => '0');
    variable r141 : std_logic_vector(0 to 0) := (others => '0');
    variable r139 : std_logic_vector(0 to 0) := (others => '0');
    variable r137 : std_logic_vector(0 to 0) := (others => '0');
    variable r135 : std_logic_vector(0 to 0) := (others => '0');
    variable r133 : std_logic_vector(0 to 0) := (others => '0');
    variable r131 : std_logic_vector(0 to 7) := (others => '0');
    variable r129 : std_logic_vector(0 to 0) := (others => '0');
    variable r127 : std_logic_vector(0 to 0) := (others => '0');
    variable r125 : std_logic_vector(0 to 0) := (others => '0');
    variable r123 : std_logic_vector(0 to 0) := (others => '0');
    variable r121 : std_logic_vector(0 to 0) := (others => '0');
    variable r119 : std_logic_vector(0 to 0) := (others => '0');
    variable r117 : std_logic_vector(0 to 0) := (others => '0');
    variable r115 : std_logic_vector(0 to 0) := (others => '0');
    variable r113 : std_logic_vector(0 to 7) := (others => '0');
    variable r111 : std_logic_vector(0 to 0) := (others => '0');
    variable r109 : std_logic_vector(0 to 0) := (others => '0');
    variable r107 : std_logic_vector(0 to 0) := (others => '0');
    variable r105 : std_logic_vector(0 to 0) := (others => '0');
    variable r103 : std_logic_vector(0 to 0) := (others => '0');
    variable r101 : std_logic_vector(0 to 0) := (others => '0');
    variable r99 : std_logic_vector(0 to 0) := (others => '0');
    variable r97 : std_logic_vector(0 to 0) := (others => '0');
    variable r95 : std_logic_vector(0 to 7) := (others => '0');
    variable r93 : std_logic_vector(0 to 0) := (others => '0');
    variable r91 : std_logic_vector(0 to 0) := (others => '0');
    variable r89 : std_logic_vector(0 to 0) := (others => '0');
    variable r87 : std_logic_vector(0 to 0) := (others => '0');
    variable r85 : std_logic_vector(0 to 0) := (others => '0');
    variable r83 : std_logic_vector(0 to 0) := (others => '0');
    variable r81 : std_logic_vector(0 to 0) := (others => '0');
    variable r79 : std_logic_vector(0 to 0) := (others => '0');
    variable r77 : std_logic_vector(0 to 7) := (others => '0');
    variable r75 : std_logic_vector(0 to 0) := (others => '0');
    variable r73 : std_logic_vector(0 to 0) := (others => '0');
    variable r71 : std_logic_vector(0 to 0) := (others => '0');
    variable r69 : std_logic_vector(0 to 0) := (others => '0');
    variable r67 : std_logic_vector(0 to 0) := (others => '0');
    variable r65 : std_logic_vector(0 to 0) := (others => '0');
    variable r63 : std_logic_vector(0 to 0) := (others => '0');
    variable r61 : std_logic_vector(0 to 0) := (others => '0');
    variable r59 : std_logic_vector(0 to 7) := (others => '0');
    variable r57 : std_logic_vector(0 to 0) := (others => '0');
    variable r55 : std_logic_vector(0 to 0) := (others => '0');
    variable r53 : std_logic_vector(0 to 0) := (others => '0');
    variable r51 : std_logic_vector(0 to 0) := (others => '0');
    variable r49 : std_logic_vector(0 to 0) := (others => '0');
    variable r47 : std_logic_vector(0 to 0) := (others => '0');
    variable r45 : std_logic_vector(0 to 0) := (others => '0');
    variable r43 : std_logic_vector(0 to 0) := (others => '0');
    variable r41 : std_logic_vector(0 to 7) := (others => '0');
    variable r39 : std_logic_vector(0 to 0) := (others => '0');
    variable r37 : std_logic_vector(0 to 0) := (others => '0');
    variable r35 : std_logic_vector(0 to 0) := (others => '0');
    variable r33 : std_logic_vector(0 to 0) := (others => '0');
    variable r31 : std_logic_vector(0 to 0) := (others => '0');
    variable r29 : std_logic_vector(0 to 0) := (others => '0');
    variable r27 : std_logic_vector(0 to 0) := (others => '0');
    variable r25 : std_logic_vector(0 to 0) := (others => '0');
    variable r23 : std_logic_vector(0 to 7) := (others => '0');
    variable r21 : std_logic_vector(0 to 0) := (others => '0');
    variable r19 : std_logic_vector(0 to 0) := (others => '0');
    variable r17 : std_logic_vector(0 to 0) := (others => '0');
    variable r15 : std_logic_vector(0 to 0) := (others => '0');
    variable r13 : std_logic_vector(0 to 0) := (others => '0');
    variable r11 : std_logic_vector(0 to 0) := (others => '0');
    variable r9 : std_logic_vector(0 to 0) := (others => '0');
    variable r7 : std_logic_vector(0 to 0) := (others => '0');
  begin
    r7 := "1";
    r9 := "1";
    r11 := "1";
    r13 := "1";
    r15 := "1";
    r17 := "1";
    r19 := "1";
    r21 := "1";
    r23 := (r7 & r9 & r11 & r13 & r15 & r17 & r19 & r21);
    r25 := "1";
    r27 := "1";
    r29 := "1";
    r31 := "1";
    r33 := "1";
    r35 := "1";
    r37 := "1";
    r39 := "1";
    r41 := (r25 & r27 & r29 & r31 & r33 & r35 & r37 & r39);
    r43 := "1";
    r45 := "1";
    r47 := "1";
    r49 := "1";
    r51 := "1";
    r53 := "1";
    r55 := "1";
    r57 := "1";
    r59 := (r43 & r45 & r47 & r49 & r51 & r53 & r55 & r57);
    r61 := "1";
    r63 := "1";
    r65 := "1";
    r67 := "1";
    r69 := "1";
    r71 := "1";
    r73 := "1";
    r75 := "1";
    r77 := (r61 & r63 & r65 & r67 & r69 & r71 & r73 & r75);
    r79 := "1";
    r81 := "1";
    r83 := "1";
    r85 := "1";
    r87 := "1";
    r89 := "1";
    r91 := "1";
    r93 := "1";
    r95 := (r79 & r81 & r83 & r85 & r87 & r89 & r91 & r93);
    r97 := "1";
    r99 := "1";
    r101 := "1";
    r103 := "1";
    r105 := "1";
    r107 := "1";
    r109 := "1";
    r111 := "1";
    r113 := (r97 & r99 & r101 & r103 & r105 & r107 & r109 & r111);
    r115 := "1";
    r117 := "1";
    r119 := "1";
    r121 := "1";
    r123 := "1";
    r125 := "1";
    r127 := "1";
    r129 := "1";
    r131 := (r115 & r117 & r119 & r121 & r123 & r125 & r127 & r129);
    r133 := "1";
    r135 := "1";
    r137 := "1";
    r139 := "1";
    r141 := "1";
    r143 := "1";
    r145 := "1";
    r147 := "1";
    r149 := (r133 & r135 & r137 & r139 & r141 & r143 & r145 & r147);
    r151 := "1";
    r153 := "1";
    r155 := "1";
    r157 := "1";
    r159 := "1";
    r161 := "1";
    r163 := "1";
    r165 := "1";
    r167 := (r151 & r153 & r155 & r157 & r159 & r161 & r163 & r165);
    r169 := "1";
    r171 := "1";
    r173 := "1";
    r175 := "1";
    r177 := "1";
    r179 := "1";
    r181 := "1";
    r183 := "1";
    r185 := (r169 & r171 & r173 & r175 & r177 & r179 & r181 & r183);
    r187 := "1";
    r189 := "1";
    r191 := "1";
    r193 := "1";
    r195 := "1";
    r197 := "1";
    r199 := "1";
    r201 := "1";
    r203 := (r187 & r189 & r191 & r193 & r195 & r197 & r199 & r201);
    r205 := "1";
    r207 := "1";
    r209 := "1";
    r211 := "1";
    r213 := "1";
    r215 := "1";
    r217 := "1";
    r219 := "1";
    r221 := (r205 & r207 & r209 & r211 & r213 & r215 & r217 & r219);
    r223 := "1";
    r225 := "1";
    r227 := "1";
    r229 := "1";
    r231 := "1";
    r233 := "1";
    r235 := "1";
    r237 := "1";
    r239 := (r223 & r225 & r227 & r229 & r231 & r233 & r235 & r237);
    r241 := "1";
    r243 := "1";
    r245 := "1";
    r247 := "1";
    r249 := "1";
    r251 := "1";
    r253 := "1";
    r255 := "1";
    r257 := (r241 & r243 & r245 & r247 & r249 & r251 & r253 & r255);
    r259 := "1";
    r261 := "1";
    r263 := "1";
    r265 := "1";
    r267 := "1";
    r269 := "1";
    r271 := "1";
    r273 := "1";
    r275 := (r259 & r261 & r263 & r265 & r267 & r269 & r271 & r273);
    r277 := "1";
    r279 := "1";
    r281 := "1";
    r283 := "1";
    r285 := "1";
    r287 := "1";
    r289 := "1";
    r291 := "1";
    r293 := (r277 & r279 & r281 & r283 & r285 & r287 & r289 & r291);
    r295 := "1";
    r297 := "1";
    r299 := "1";
    r301 := "1";
    r303 := "1";
    r305 := "1";
    r307 := "1";
    r309 := "1";
    r311 := (r295 & r297 & r299 & r301 & r303 & r305 & r307 & r309);
    r313 := "1";
    r315 := "1";
    r317 := "1";
    r319 := "1";
    r321 := "1";
    r323 := "1";
    r325 := "1";
    r327 := "1";
    r329 := (r313 & r315 & r317 & r319 & r321 & r323 & r325 & r327);
    r331 := "1";
    r333 := "1";
    r335 := "1";
    r337 := "1";
    r339 := "1";
    r341 := "1";
    r343 := "1";
    r345 := "1";
    r347 := (r331 & r333 & r335 & r337 & r339 & r341 & r343 & r345);
    r349 := "1";
    r351 := "1";
    r353 := "1";
    r355 := "1";
    r357 := "1";
    r359 := "1";
    r361 := "1";
    r363 := "1";
    r365 := (r349 & r351 & r353 & r355 & r357 & r359 & r361 & r363);
    r367 := "1";
    r369 := "1";
    r371 := "1";
    r373 := "1";
    r375 := "1";
    r377 := "1";
    r379 := "1";
    r381 := "1";
    r383 := (r367 & r369 & r371 & r373 & r375 & r377 & r379 & r381);
    r385 := "1";
    r387 := "1";
    r389 := "1";
    r391 := "1";
    r393 := "1";
    r395 := "1";
    r397 := "1";
    r399 := "1";
    r401 := (r385 & r387 & r389 & r391 & r393 & r395 & r397 & r399);
    r403 := "1";
    r405 := "1";
    r407 := "1";
    r409 := "1";
    r411 := "1";
    r413 := "1";
    r415 := "1";
    r417 := "1";
    r419 := (r403 & r405 & r407 & r409 & r411 & r413 & r415 & r417);
    r421 := "1";
    r423 := "1";
    r425 := "1";
    r427 := "1";
    r429 := "1";
    r431 := "1";
    r433 := "1";
    r435 := "1";
    r437 := (r421 & r423 & r425 & r427 & r429 & r431 & r433 & r435);
    r439 := "1";
    r441 := "1";
    r443 := "1";
    r445 := "1";
    r447 := "1";
    r449 := "1";
    r451 := "1";
    r453 := "1";
    r455 := (r439 & r441 & r443 & r445 & r447 & r449 & r451 & r453);
    r457 := "1";
    r459 := "1";
    r461 := "1";
    r463 := "1";
    r465 := "1";
    r467 := "1";
    r469 := "1";
    r471 := "1";
    r473 := (r457 & r459 & r461 & r463 & r465 & r467 & r469 & r471);
    r475 := "1";
    r477 := "1";
    r479 := "1";
    r481 := "1";
    r483 := "1";
    r485 := "1";
    r487 := "1";
    r489 := "1";
    r491 := (r475 & r477 & r479 & r481 & r483 & r485 & r487 & r489);
    r493 := "1";
    r495 := "1";
    r497 := "1";
    r499 := "1";
    r501 := "1";
    r503 := "1";
    r505 := "1";
    r507 := "1";
    r509 := (r493 & r495 & r497 & r499 & r501 & r503 & r505 & r507);
    r511 := "1";
    r513 := "1";
    r515 := "1";
    r517 := "1";
    r519 := "1";
    r521 := "1";
    r523 := "1";
    r525 := "1";
    r527 := (r511 & r513 & r515 & r517 & r519 & r521 & r523 & r525);
    r529 := "1";
    r531 := "1";
    r533 := "1";
    r535 := "1";
    r537 := "1";
    r539 := "1";
    r541 := "1";
    r543 := "1";
    r545 := (r529 & r531 & r533 & r535 & r537 & r539 & r541 & r543);
    r547 := "1";
    r549 := "1";
    r551 := "1";
    r553 := "1";
    r555 := "1";
    r557 := "1";
    r559 := "1";
    r561 := "1";
    r563 := (r547 & r549 & r551 & r553 & r555 & r557 & r559 & r561);
    r565 := "1";
    r567 := "1";
    r569 := "1";
    r571 := "1";
    r573 := "1";
    r575 := "1";
    r577 := "1";
    r579 := "1";
    r581 := (r565 & r567 & r569 & r571 & r573 & r575 & r577 & r579);
    r583 := "1";
    r585 := "1";
    r587 := "1";
    r589 := "1";
    r591 := "1";
    r593 := "1";
    r595 := "1";
    r597 := "1";
    r599 := (r583 & r585 & r587 & r589 & r591 & r593 & r595 & r597);
    r601 := "1";
    r603 := "1";
    r605 := "1";
    r607 := "1";
    r609 := "1";
    r611 := "1";
    r613 := "1";
    r615 := "1";
    r617 := (r601 & r603 & r605 & r607 & r609 & r611 & r613 & r615);
    r619 := "1";
    r621 := "1";
    r623 := "1";
    r625 := "1";
    r627 := "1";
    r629 := "1";
    r631 := "1";
    r633 := "1";
    r635 := (r619 & r621 & r623 & r625 & r627 & r629 & r631 & r633);
    r637 := "1";
    r639 := "1";
    r641 := "1";
    r643 := "1";
    r645 := "1";
    r647 := "1";
    r649 := "1";
    r651 := "1";
    r653 := (r637 & r639 & r641 & r643 & r645 & r647 & r649 & r651);
    r655 := "1";
    r657 := "1";
    r659 := "1";
    r661 := "1";
    r663 := "1";
    r665 := "1";
    r667 := "1";
    r669 := "1";
    r671 := (r655 & r657 & r659 & r661 & r663 & r665 & r667 & r669);
    r673 := "1";
    r675 := "1";
    r677 := "1";
    r679 := "1";
    r681 := "1";
    r683 := "1";
    r685 := "1";
    r687 := "1";
    r689 := (r673 & r675 & r677 & r679 & r681 & r683 & r685 & r687);
    r691 := "1";
    r693 := "1";
    r695 := "1";
    r697 := "1";
    r699 := "1";
    r701 := "1";
    r703 := "1";
    r705 := "1";
    r707 := (r691 & r693 & r695 & r697 & r699 & r701 & r703 & r705);
    r709 := "1";
    r711 := "1";
    r713 := "1";
    r715 := "1";
    r717 := "1";
    r719 := "1";
    r721 := "1";
    r723 := "1";
    r725 := (r709 & r711 & r713 & r715 & r717 & r719 & r721 & r723);
    r727 := "1";
    r729 := "1";
    r731 := "1";
    r733 := "1";
    r735 := "1";
    r737 := "1";
    r739 := "1";
    r741 := "1";
    r743 := (r727 & r729 & r731 & r733 & r735 & r737 & r739 & r741);
    r745 := "1";
    r747 := "1";
    r749 := "1";
    r751 := "1";
    r753 := "1";
    r755 := "1";
    r757 := "1";
    r759 := "1";
    r761 := (r745 & r747 & r749 & r751 & r753 & r755 & r757 & r759);
    r763 := "1";
    r765 := "1";
    r767 := "1";
    r769 := "1";
    r771 := "1";
    r773 := "1";
    r775 := "1";
    r777 := "1";
    r779 := (r763 & r765 & r767 & r769 & r771 & r773 & r775 & r777);
    r781 := "1";
    r783 := "1";
    r785 := "1";
    r787 := "1";
    r789 := "1";
    r791 := "1";
    r793 := "1";
    r795 := "1";
    r797 := (r781 & r783 & r785 & r787 & r789 & r791 & r793 & r795);
    r799 := "1";
    r801 := "1";
    r803 := "1";
    r805 := "1";
    r807 := "1";
    r809 := "1";
    r811 := "1";
    r813 := "1";
    r815 := (r799 & r801 & r803 & r805 & r807 & r809 & r811 & r813);
    r817 := "1";
    r819 := "1";
    r821 := "1";
    r823 := "1";
    r825 := "1";
    r827 := "1";
    r829 := "1";
    r831 := "1";
    r833 := (r817 & r819 & r821 & r823 & r825 & r827 & r829 & r831);
    r835 := "1";
    r837 := "1";
    r839 := "1";
    r841 := "1";
    r843 := "1";
    r845 := "1";
    r847 := "1";
    r849 := "1";
    r851 := (r835 & r837 & r839 & r841 & r843 & r845 & r847 & r849);
    r853 := "1";
    r855 := "1";
    r857 := "1";
    r859 := "1";
    r861 := "1";
    r863 := "1";
    r865 := "1";
    r867 := "1";
    r869 := (r853 & r855 & r857 & r859 & r861 & r863 & r865 & r867);
    r871 := "1";
    r873 := "1";
    r875 := "1";
    r877 := "1";
    r879 := "1";
    r881 := "1";
    r883 := "1";
    r885 := "1";
    r887 := (r871 & r873 & r875 & r877 & r879 & r881 & r883 & r885);
    r889 := "1";
    r891 := "1";
    r893 := "1";
    r895 := "1";
    r897 := "1";
    r899 := "1";
    r901 := "1";
    r903 := "1";
    r905 := (r889 & r891 & r893 & r895 & r897 & r899 & r901 & r903);
    r907 := "1";
    r909 := "1";
    r911 := "1";
    r913 := "1";
    r915 := "1";
    r917 := "1";
    r919 := "1";
    r921 := "1";
    r923 := (r907 & r909 & r911 & r913 & r915 & r917 & r919 & r921);
    r925 := "1";
    r927 := "1";
    r929 := "1";
    r931 := "1";
    r933 := "1";
    r935 := "1";
    r937 := "1";
    r939 := "1";
    r941 := (r925 & r927 & r929 & r931 & r933 & r935 & r937 & r939);
    r943 := "1";
    r945 := "1";
    r947 := "1";
    r949 := "1";
    r951 := "1";
    r953 := "1";
    r955 := "1";
    r957 := "1";
    r959 := (r943 & r945 & r947 & r949 & r951 & r953 & r955 & r957);
    r961 := "1";
    r963 := "1";
    r965 := "1";
    r967 := "1";
    r969 := "1";
    r971 := "1";
    r973 := "1";
    r975 := "1";
    r977 := (r961 & r963 & r965 & r967 & r969 & r971 & r973 & r975);
    r979 := "1";
    r981 := "1";
    r983 := "1";
    r985 := "1";
    r987 := "1";
    r989 := "1";
    r991 := "1";
    r993 := "1";
    r995 := (r979 & r981 & r983 & r985 & r987 & r989 & r991 & r993);
    r997 := "1";
    r999 := "1";
    r1001 := "1";
    r1003 := "1";
    r1005 := "1";
    r1007 := "1";
    r1009 := "1";
    r1011 := "1";
    r1013 := (r997 & r999 & r1001 & r1003 & r1005 & r1007 & r1009 & r1011);
    r1015 := "1";
    r1017 := "1";
    r1019 := "1";
    r1021 := "1";
    r1023 := "1";
    r1025 := "1";
    r1027 := "1";
    r1029 := "1";
    r1031 := (r1015 & r1017 & r1019 & r1021 & r1023 & r1025 & r1027 & r1029);
    r1033 := "1";
    r1035 := "1";
    r1037 := "1";
    r1039 := "1";
    r1041 := "1";
    r1043 := "1";
    r1045 := "1";
    r1047 := "1";
    r1049 := (r1033 & r1035 & r1037 & r1039 & r1041 & r1043 & r1045 & r1047);
    r1051 := "1";
    r1053 := "1";
    r1055 := "1";
    r1057 := "1";
    r1059 := "1";
    r1061 := "1";
    r1063 := "1";
    r1065 := "1";
    r1067 := (r1051 & r1053 & r1055 & r1057 & r1059 & r1061 & r1063 & r1065);
    r1069 := "1";
    r1071 := "1";
    r1073 := "1";
    r1075 := "1";
    r1077 := "1";
    r1079 := "1";
    r1081 := "1";
    r1083 := "1";
    r1085 := (r1069 & r1071 & r1073 & r1075 & r1077 & r1079 & r1081 & r1083);
    r1087 := "1";
    r1089 := "1";
    r1091 := "1";
    r1093 := "1";
    r1095 := "1";
    r1097 := "1";
    r1099 := "1";
    r1101 := "1";
    r1103 := (r1087 & r1089 & r1091 & r1093 & r1095 & r1097 & r1099 & r1101);
    r1105 := "1";
    r1107 := "1";
    r1109 := "1";
    r1111 := "1";
    r1113 := "1";
    r1115 := "1";
    r1117 := "1";
    r1119 := "1";
    r1121 := (r1105 & r1107 & r1109 & r1111 & r1113 & r1115 & r1117 & r1119);
    r1123 := "1";
    r1125 := "1";
    r1127 := "1";
    r1129 := "1";
    r1131 := "1";
    r1133 := "1";
    r1135 := "1";
    r1137 := "1";
    r1139 := (r1123 & r1125 & r1127 & r1129 & r1131 & r1133 & r1135 & r1137);
    r1141 := "1";
    r1143 := "1";
    r1145 := "1";
    r1147 := "1";
    r1149 := "1";
    r1151 := "1";
    r1153 := "1";
    r1155 := "1";
    r1157 := (r1141 & r1143 & r1145 & r1147 & r1149 & r1151 & r1153 & r1155);
    r1158 := (r23 & r41 & r59 & r77 & r95 & r113 & r131 & r149 & r167 & r185 & r203 & r221 & r239 & r257 & r275 & r293 & r311 & r329 & r347 & r365 & r383 & r401 & r419 & r437 & r455 & r473 & r491 & r509 & r527 & r545 & r563 & r581 & r599 & r617 & r635 & r653 & r671 & r689 & r707 & r725 & r743 & r761 & r779 & r797 & r815 & r833 & r851 & r869 & r887 & r905 & r923 & r941 & r959 & r977 & r995 & r1013 & r1031 & r1049 & r1067 & r1085 & r1103 & r1121 & r1139 & r1157);
    return r1158;
  end rewire_zerothoutput_3;

begin
  process (clk)
    variable goto_L3543 : boolean := false;
    variable goto_L3537 : boolean := false;
    variable goto_L1163 : boolean := false;
    variable goto_L1165 : boolean := false;
    variable goto_L0 : boolean := false;
    variable goto_L3544 : boolean := false;
    variable r3536 : std_logic_vector(0 to 639) := (others => '0');
    variable r3533 : std_logic_vector(0 to 511) := (others => '0');
    variable r3529 : std_logic_vector(0 to 511) := (others => '0');
    variable r3525 : std_logic_vector(0 to 127) := (others => '0');
    variable r3234 : std_logic_vector(0 to 127) := (others => '0');
    variable r3231 : std_logic_vector(0 to 127) := (others => '0');
    variable r2940 : std_logic_vector(0 to 127) := (others => '0');
    variable r1187 : std_logic_vector(0 to 511) := (others => '0');
    variable r1186 : std_logic_vector(0 to 63) := (others => '0');
    variable r1185 : std_logic_vector(0 to 63) := (others => '0');
    variable r1184 : std_logic_vector(0 to 127) := (others => '0');
    variable r1183 : std_logic_vector(0 to 127) := (others => '0');
    variable b1180 : boolean := false;
    variable b1178 : boolean := false;
    variable b1176 : boolean := false;
    variable r1174 : std_logic_vector(0 to 511) := (others => '0');
    variable r1172 : std_logic_vector(0 to 63) := (others => '0');
    variable r1170 : std_logic_vector(0 to 63) := (others => '0');
    variable r1164 : std_logic_vector(0 to 639) := (others => '0');
    variable r1162 : std_logic_vector(0 to 639) := (others => '0');
    variable r1159 : std_logic_vector(0 to 511) := (others => '0');
    variable r4 : std_logic_vector(0 to 511) := (others => '0');
    variable state : control_state := STATE0;
  begin
    if clk'event and clk='1' then
      goto_L3543 := false;
      goto_L3537 := false;
      goto_L1163 := false;
      goto_L1165 := false;
      goto_L0 := false;
      goto_L3544 := false;
      null; -- label L3543
      -- ENTER
      goto_L0 := (state = STATE0);
      if (NOT goto_L0) then
        goto_L1163 := (state = STATE1163);
        if (NOT goto_L1163) then
          goto_L3537 := (state = STATE3537);
          null; -- label L3537
          r3536 := input;
          -- got r@IU in r3536
          r1164 := r3536;
          goto_L1165 := true;
        end if;
        goto_L1165 := goto_L1165;
        if (NOT goto_L1165) then
          null; -- label L1163
          r1162 := input;
          -- got r@IV in r1162
          r1164 := r1162;
          goto_L1165 := true;
        end if;
        goto_L1165 := goto_L1165;
        null; -- label L1165
        -- step in
        -- got x@IP in r1164
        -- final pat
        r1170 := r1164(0 to 63);
        r1172 := r1164(64 to 127);
        r1174 := r1164(128 to 639);
        b1176 := true;
        b1178 := true;
        b1180 := true;
        r3231 := rewire_key1_2939;
        r3525 := rewire_key2_3233;
        -- got b0@IQ in r1170
        -- got b1@IR in r1172
        r3529 := rewire_buildSalsa256_1182(r3231,r3525,r1170,r1172);
        -- got y@IT in r3529
        -- got b64@IS in r1174
        r3533 := xor512(r3529,r1174);
        output <= r3533;
        state := STATE3537;
        goto_L3544 := true;
      end if;
      goto_L3544 := goto_L3544;
      if (NOT goto_L3544) then
        null; -- label L0
        -- START
        -- foo in
        r1159 := rewire_zerothoutput_3;
        output <= r1159;
        state := STATE1163;
        goto_L3544 := true;
      end if;
      goto_L3544 := goto_L3544;
      null; -- label L3544
      -- EXIT
    end if;
  end process;
end behavioral;
library ieee;
use ieee.std_logic_1164.all;
-- Uncomment the following line if VHDL primitives are in use.
-- use prims.all;
entity main is
  Port ( clk : in std_logic ;
         input : in std_logic_vector (0 to 639);
         output : out std_logic_vector (0 to 511));
end main;
architecture structural of main is
begin
  dev : entity work.rwcomp0(behavioral)
    port map (clk,input,output);
    

end structural;
