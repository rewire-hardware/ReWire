library ieee;
use ieee.std_logic_1164.all;
-- Uncomment the following line if VHDL primitives are in use.
use work.prims.all;
entity rwcomp0 is
  Port ( clk : in std_logic ;
         input : in std_logic_vector (0 to 127);
         output : out std_logic_vector (0 to 511));
end rwcomp0;

architecture behavioral of rwcomp0 is
  type control_state is (STATE0,STATE1163,STATE3530);
  function rewire_key2_3229 return std_logic_vector;
  function rewire_key1_2935 return std_logic_vector;
  function rewire_buildSalsa256_1178(r1179 : std_logic_vector ; r1180 : std_logic_vector ; r1181 : std_logic_vector ; r1182 : std_logic_vector) return std_logic_vector;
  function rewire_salsaHash_1654(r1655 : std_logic_vector) return std_logic_vector;
  function rewire_impwords_2598(r2599 : std_logic_vector) return std_logic_vector;
  function rewire_littleendian_2732(r2733 : std_logic_vector) return std_logic_vector;
  function rewire_w8to16le_2827(r2828 : std_logic_vector ; r2829 : std_logic_vector) return std_logic_vector;
  function rewire_w16tow32le_2746(r2747 : std_logic_vector ; r2748 : std_logic_vector) return std_logic_vector;
  function rewire_salsaHashp_1974(r1975 : std_logic_vector) return std_logic_vector;
  function rewire_doubleRound_2012(r2013 : std_logic_vector) return std_logic_vector;
  function rewire_columnRound_2432(r2433 : std_logic_vector) return std_logic_vector;
  function rewire_rowRound_2015(r2016 : std_logic_vector) return std_logic_vector;
  function rewire_quarterRound_2053(r2054 : std_logic_vector) return std_logic_vector;
  function rewire_rot18_2292(r2293 : std_logic_vector) return std_logic_vector;
  function rewire_rot13_2217(r2218 : std_logic_vector) return std_logic_vector;
  function rewire_rot9_2142(r2143 : std_logic_vector) return std_logic_vector;
  function rewire_rot7_2067(r2068 : std_logic_vector) return std_logic_vector;
  function rewire_expwords_1657(r1658 : std_logic_vector) return std_logic_vector;
  function rewire_littleendianp_1695(r1696 : std_logic_vector) return std_logic_vector;
  function rewire_sigma3_1529 return std_logic_vector;
  function rewire_sigma2_1452 return std_logic_vector;
  function rewire_sigma1_1375 return std_logic_vector;
  function rewire_sigma0_1298 return std_logic_vector;
  function rewire_zerothoutput_3 return std_logic_vector;

  function rewire_key2_3229 return std_logic_vector
  is
    variable r3520 : std_logic_vector(0 to 127) := (others => '0');
    variable r3519 : std_logic_vector(0 to 7) := (others => '0');
    variable r3517 : std_logic_vector(0 to 0) := (others => '0');
    variable r3515 : std_logic_vector(0 to 0) := (others => '0');
    variable r3513 : std_logic_vector(0 to 0) := (others => '0');
    variable r3511 : std_logic_vector(0 to 0) := (others => '0');
    variable r3509 : std_logic_vector(0 to 0) := (others => '0');
    variable r3507 : std_logic_vector(0 to 0) := (others => '0');
    variable r3505 : std_logic_vector(0 to 0) := (others => '0');
    variable r3503 : std_logic_vector(0 to 0) := (others => '0');
    variable r3501 : std_logic_vector(0 to 7) := (others => '0');
    variable r3499 : std_logic_vector(0 to 0) := (others => '0');
    variable r3497 : std_logic_vector(0 to 0) := (others => '0');
    variable r3495 : std_logic_vector(0 to 0) := (others => '0');
    variable r3493 : std_logic_vector(0 to 0) := (others => '0');
    variable r3491 : std_logic_vector(0 to 0) := (others => '0');
    variable r3489 : std_logic_vector(0 to 0) := (others => '0');
    variable r3487 : std_logic_vector(0 to 0) := (others => '0');
    variable r3485 : std_logic_vector(0 to 0) := (others => '0');
    variable r3483 : std_logic_vector(0 to 7) := (others => '0');
    variable r3481 : std_logic_vector(0 to 0) := (others => '0');
    variable r3479 : std_logic_vector(0 to 0) := (others => '0');
    variable r3477 : std_logic_vector(0 to 0) := (others => '0');
    variable r3475 : std_logic_vector(0 to 0) := (others => '0');
    variable r3473 : std_logic_vector(0 to 0) := (others => '0');
    variable r3471 : std_logic_vector(0 to 0) := (others => '0');
    variable r3469 : std_logic_vector(0 to 0) := (others => '0');
    variable r3467 : std_logic_vector(0 to 0) := (others => '0');
    variable r3465 : std_logic_vector(0 to 7) := (others => '0');
    variable r3463 : std_logic_vector(0 to 0) := (others => '0');
    variable r3461 : std_logic_vector(0 to 0) := (others => '0');
    variable r3459 : std_logic_vector(0 to 0) := (others => '0');
    variable r3457 : std_logic_vector(0 to 0) := (others => '0');
    variable r3455 : std_logic_vector(0 to 0) := (others => '0');
    variable r3453 : std_logic_vector(0 to 0) := (others => '0');
    variable r3451 : std_logic_vector(0 to 0) := (others => '0');
    variable r3449 : std_logic_vector(0 to 0) := (others => '0');
    variable r3447 : std_logic_vector(0 to 7) := (others => '0');
    variable r3445 : std_logic_vector(0 to 0) := (others => '0');
    variable r3443 : std_logic_vector(0 to 0) := (others => '0');
    variable r3441 : std_logic_vector(0 to 0) := (others => '0');
    variable r3439 : std_logic_vector(0 to 0) := (others => '0');
    variable r3437 : std_logic_vector(0 to 0) := (others => '0');
    variable r3435 : std_logic_vector(0 to 0) := (others => '0');
    variable r3433 : std_logic_vector(0 to 0) := (others => '0');
    variable r3431 : std_logic_vector(0 to 0) := (others => '0');
    variable r3429 : std_logic_vector(0 to 7) := (others => '0');
    variable r3427 : std_logic_vector(0 to 0) := (others => '0');
    variable r3425 : std_logic_vector(0 to 0) := (others => '0');
    variable r3423 : std_logic_vector(0 to 0) := (others => '0');
    variable r3421 : std_logic_vector(0 to 0) := (others => '0');
    variable r3419 : std_logic_vector(0 to 0) := (others => '0');
    variable r3417 : std_logic_vector(0 to 0) := (others => '0');
    variable r3415 : std_logic_vector(0 to 0) := (others => '0');
    variable r3413 : std_logic_vector(0 to 0) := (others => '0');
    variable r3411 : std_logic_vector(0 to 7) := (others => '0');
    variable r3409 : std_logic_vector(0 to 0) := (others => '0');
    variable r3407 : std_logic_vector(0 to 0) := (others => '0');
    variable r3405 : std_logic_vector(0 to 0) := (others => '0');
    variable r3403 : std_logic_vector(0 to 0) := (others => '0');
    variable r3401 : std_logic_vector(0 to 0) := (others => '0');
    variable r3399 : std_logic_vector(0 to 0) := (others => '0');
    variable r3397 : std_logic_vector(0 to 0) := (others => '0');
    variable r3395 : std_logic_vector(0 to 0) := (others => '0');
    variable r3393 : std_logic_vector(0 to 7) := (others => '0');
    variable r3391 : std_logic_vector(0 to 0) := (others => '0');
    variable r3389 : std_logic_vector(0 to 0) := (others => '0');
    variable r3387 : std_logic_vector(0 to 0) := (others => '0');
    variable r3385 : std_logic_vector(0 to 0) := (others => '0');
    variable r3383 : std_logic_vector(0 to 0) := (others => '0');
    variable r3381 : std_logic_vector(0 to 0) := (others => '0');
    variable r3379 : std_logic_vector(0 to 0) := (others => '0');
    variable r3377 : std_logic_vector(0 to 0) := (others => '0');
    variable r3375 : std_logic_vector(0 to 7) := (others => '0');
    variable r3373 : std_logic_vector(0 to 0) := (others => '0');
    variable r3371 : std_logic_vector(0 to 0) := (others => '0');
    variable r3369 : std_logic_vector(0 to 0) := (others => '0');
    variable r3367 : std_logic_vector(0 to 0) := (others => '0');
    variable r3365 : std_logic_vector(0 to 0) := (others => '0');
    variable r3363 : std_logic_vector(0 to 0) := (others => '0');
    variable r3361 : std_logic_vector(0 to 0) := (others => '0');
    variable r3359 : std_logic_vector(0 to 0) := (others => '0');
    variable r3357 : std_logic_vector(0 to 7) := (others => '0');
    variable r3355 : std_logic_vector(0 to 0) := (others => '0');
    variable r3353 : std_logic_vector(0 to 0) := (others => '0');
    variable r3351 : std_logic_vector(0 to 0) := (others => '0');
    variable r3349 : std_logic_vector(0 to 0) := (others => '0');
    variable r3347 : std_logic_vector(0 to 0) := (others => '0');
    variable r3345 : std_logic_vector(0 to 0) := (others => '0');
    variable r3343 : std_logic_vector(0 to 0) := (others => '0');
    variable r3341 : std_logic_vector(0 to 0) := (others => '0');
    variable r3339 : std_logic_vector(0 to 7) := (others => '0');
    variable r3337 : std_logic_vector(0 to 0) := (others => '0');
    variable r3335 : std_logic_vector(0 to 0) := (others => '0');
    variable r3333 : std_logic_vector(0 to 0) := (others => '0');
    variable r3331 : std_logic_vector(0 to 0) := (others => '0');
    variable r3329 : std_logic_vector(0 to 0) := (others => '0');
    variable r3327 : std_logic_vector(0 to 0) := (others => '0');
    variable r3325 : std_logic_vector(0 to 0) := (others => '0');
    variable r3323 : std_logic_vector(0 to 0) := (others => '0');
    variable r3321 : std_logic_vector(0 to 7) := (others => '0');
    variable r3319 : std_logic_vector(0 to 0) := (others => '0');
    variable r3317 : std_logic_vector(0 to 0) := (others => '0');
    variable r3315 : std_logic_vector(0 to 0) := (others => '0');
    variable r3313 : std_logic_vector(0 to 0) := (others => '0');
    variable r3311 : std_logic_vector(0 to 0) := (others => '0');
    variable r3309 : std_logic_vector(0 to 0) := (others => '0');
    variable r3307 : std_logic_vector(0 to 0) := (others => '0');
    variable r3305 : std_logic_vector(0 to 0) := (others => '0');
    variable r3303 : std_logic_vector(0 to 7) := (others => '0');
    variable r3301 : std_logic_vector(0 to 0) := (others => '0');
    variable r3299 : std_logic_vector(0 to 0) := (others => '0');
    variable r3297 : std_logic_vector(0 to 0) := (others => '0');
    variable r3295 : std_logic_vector(0 to 0) := (others => '0');
    variable r3293 : std_logic_vector(0 to 0) := (others => '0');
    variable r3291 : std_logic_vector(0 to 0) := (others => '0');
    variable r3289 : std_logic_vector(0 to 0) := (others => '0');
    variable r3287 : std_logic_vector(0 to 0) := (others => '0');
    variable r3285 : std_logic_vector(0 to 7) := (others => '0');
    variable r3283 : std_logic_vector(0 to 0) := (others => '0');
    variable r3281 : std_logic_vector(0 to 0) := (others => '0');
    variable r3279 : std_logic_vector(0 to 0) := (others => '0');
    variable r3277 : std_logic_vector(0 to 0) := (others => '0');
    variable r3275 : std_logic_vector(0 to 0) := (others => '0');
    variable r3273 : std_logic_vector(0 to 0) := (others => '0');
    variable r3271 : std_logic_vector(0 to 0) := (others => '0');
    variable r3269 : std_logic_vector(0 to 0) := (others => '0');
    variable r3267 : std_logic_vector(0 to 7) := (others => '0');
    variable r3265 : std_logic_vector(0 to 0) := (others => '0');
    variable r3263 : std_logic_vector(0 to 0) := (others => '0');
    variable r3261 : std_logic_vector(0 to 0) := (others => '0');
    variable r3259 : std_logic_vector(0 to 0) := (others => '0');
    variable r3257 : std_logic_vector(0 to 0) := (others => '0');
    variable r3255 : std_logic_vector(0 to 0) := (others => '0');
    variable r3253 : std_logic_vector(0 to 0) := (others => '0');
    variable r3251 : std_logic_vector(0 to 0) := (others => '0');
    variable r3249 : std_logic_vector(0 to 7) := (others => '0');
    variable r3247 : std_logic_vector(0 to 0) := (others => '0');
    variable r3245 : std_logic_vector(0 to 0) := (others => '0');
    variable r3243 : std_logic_vector(0 to 0) := (others => '0');
    variable r3241 : std_logic_vector(0 to 0) := (others => '0');
    variable r3239 : std_logic_vector(0 to 0) := (others => '0');
    variable r3237 : std_logic_vector(0 to 0) := (others => '0');
    variable r3235 : std_logic_vector(0 to 0) := (others => '0');
    variable r3233 : std_logic_vector(0 to 0) := (others => '0');
    variable EMPTY : std_logic_vector(0 to -1) := (others => '0');
  begin
    r3233 := "1";
    r3235 := "0";
    r3237 := "0";
    r3239 := "0";
    r3241 := "1";
    r3243 := "0";
    r3245 := "0";
    r3247 := "0";
    r3249 := (r3233 & r3235 & r3237 & r3239 & r3241 & r3243 & r3245 & r3247);
    r3251 := "0";
    r3253 := "1";
    r3255 := "0";
    r3257 := "0";
    r3259 := "1";
    r3261 := "0";
    r3263 := "0";
    r3265 := "0";
    r3267 := (r3251 & r3253 & r3255 & r3257 & r3259 & r3261 & r3263 & r3265);
    r3269 := "1";
    r3271 := "1";
    r3273 := "0";
    r3275 := "0";
    r3277 := "1";
    r3279 := "0";
    r3281 := "0";
    r3283 := "0";
    r3285 := (r3269 & r3271 & r3273 & r3275 & r3277 & r3279 & r3281 & r3283);
    r3287 := "0";
    r3289 := "0";
    r3291 := "1";
    r3293 := "0";
    r3295 := "1";
    r3297 := "0";
    r3299 := "0";
    r3301 := "0";
    r3303 := (r3287 & r3289 & r3291 & r3293 & r3295 & r3297 & r3299 & r3301);
    r3305 := "1";
    r3307 := "0";
    r3309 := "1";
    r3311 := "0";
    r3313 := "1";
    r3315 := "0";
    r3317 := "0";
    r3319 := "0";
    r3321 := (r3305 & r3307 & r3309 & r3311 & r3313 & r3315 & r3317 & r3319);
    r3323 := "0";
    r3325 := "1";
    r3327 := "1";
    r3329 := "0";
    r3331 := "1";
    r3333 := "0";
    r3335 := "0";
    r3337 := "0";
    r3339 := (r3323 & r3325 & r3327 & r3329 & r3331 & r3333 & r3335 & r3337);
    r3341 := "1";
    r3343 := "1";
    r3345 := "1";
    r3347 := "0";
    r3349 := "1";
    r3351 := "0";
    r3353 := "0";
    r3355 := "0";
    r3357 := (r3341 & r3343 & r3345 & r3347 & r3349 & r3351 & r3353 & r3355);
    r3359 := "0";
    r3361 := "0";
    r3363 := "0";
    r3365 := "1";
    r3367 := "1";
    r3369 := "0";
    r3371 := "0";
    r3373 := "0";
    r3375 := (r3359 & r3361 & r3363 & r3365 & r3367 & r3369 & r3371 & r3373);
    r3377 := "1";
    r3379 := "0";
    r3381 := "0";
    r3383 := "1";
    r3385 := "1";
    r3387 := "0";
    r3389 := "0";
    r3391 := "0";
    r3393 := (r3377 & r3379 & r3381 & r3383 & r3385 & r3387 & r3389 & r3391);
    r3395 := "0";
    r3397 := "1";
    r3399 := "0";
    r3401 := "1";
    r3403 := "1";
    r3405 := "0";
    r3407 := "0";
    r3409 := "0";
    r3411 := (r3395 & r3397 & r3399 & r3401 & r3403 & r3405 & r3407 & r3409);
    r3413 := "1";
    r3415 := "1";
    r3417 := "0";
    r3419 := "1";
    r3421 := "1";
    r3423 := "0";
    r3425 := "0";
    r3427 := "0";
    r3429 := (r3413 & r3415 & r3417 & r3419 & r3421 & r3423 & r3425 & r3427);
    r3431 := "0";
    r3433 := "0";
    r3435 := "1";
    r3437 := "1";
    r3439 := "1";
    r3441 := "0";
    r3443 := "0";
    r3445 := "0";
    r3447 := (r3431 & r3433 & r3435 & r3437 & r3439 & r3441 & r3443 & r3445);
    r3449 := "1";
    r3451 := "0";
    r3453 := "1";
    r3455 := "1";
    r3457 := "1";
    r3459 := "0";
    r3461 := "0";
    r3463 := "0";
    r3465 := (r3449 & r3451 & r3453 & r3455 & r3457 & r3459 & r3461 & r3463);
    r3467 := "0";
    r3469 := "1";
    r3471 := "1";
    r3473 := "1";
    r3475 := "1";
    r3477 := "0";
    r3479 := "0";
    r3481 := "0";
    r3483 := (r3467 & r3469 & r3471 & r3473 & r3475 & r3477 & r3479 & r3481);
    r3485 := "1";
    r3487 := "1";
    r3489 := "1";
    r3491 := "1";
    r3493 := "1";
    r3495 := "0";
    r3497 := "0";
    r3499 := "0";
    r3501 := (r3485 & r3487 & r3489 & r3491 & r3493 & r3495 & r3497 & r3499);
    r3503 := "0";
    r3505 := "0";
    r3507 := "0";
    r3509 := "0";
    r3511 := "0";
    r3513 := "1";
    r3515 := "0";
    r3517 := "0";
    r3519 := (r3503 & r3505 & r3507 & r3509 & r3511 & r3513 & r3515 & r3517);
    r3520 := (r3249 & r3267 & r3285 & r3303 & r3321 & r3339 & r3357 & r3375 & r3393 & r3411 & r3429 & r3447 & r3465 & r3483 & r3501 & r3519);
    return r3520;
  end rewire_key2_3229;
  function rewire_key1_2935 return std_logic_vector
  is
    variable r3226 : std_logic_vector(0 to 127) := (others => '0');
    variable r3225 : std_logic_vector(0 to 7) := (others => '0');
    variable r3223 : std_logic_vector(0 to 0) := (others => '0');
    variable r3221 : std_logic_vector(0 to 0) := (others => '0');
    variable r3219 : std_logic_vector(0 to 0) := (others => '0');
    variable r3217 : std_logic_vector(0 to 0) := (others => '0');
    variable r3215 : std_logic_vector(0 to 0) := (others => '0');
    variable r3213 : std_logic_vector(0 to 0) := (others => '0');
    variable r3211 : std_logic_vector(0 to 0) := (others => '0');
    variable r3209 : std_logic_vector(0 to 0) := (others => '0');
    variable r3207 : std_logic_vector(0 to 7) := (others => '0');
    variable r3205 : std_logic_vector(0 to 0) := (others => '0');
    variable r3203 : std_logic_vector(0 to 0) := (others => '0');
    variable r3201 : std_logic_vector(0 to 0) := (others => '0');
    variable r3199 : std_logic_vector(0 to 0) := (others => '0');
    variable r3197 : std_logic_vector(0 to 0) := (others => '0');
    variable r3195 : std_logic_vector(0 to 0) := (others => '0');
    variable r3193 : std_logic_vector(0 to 0) := (others => '0');
    variable r3191 : std_logic_vector(0 to 0) := (others => '0');
    variable r3189 : std_logic_vector(0 to 7) := (others => '0');
    variable r3187 : std_logic_vector(0 to 0) := (others => '0');
    variable r3185 : std_logic_vector(0 to 0) := (others => '0');
    variable r3183 : std_logic_vector(0 to 0) := (others => '0');
    variable r3181 : std_logic_vector(0 to 0) := (others => '0');
    variable r3179 : std_logic_vector(0 to 0) := (others => '0');
    variable r3177 : std_logic_vector(0 to 0) := (others => '0');
    variable r3175 : std_logic_vector(0 to 0) := (others => '0');
    variable r3173 : std_logic_vector(0 to 0) := (others => '0');
    variable r3171 : std_logic_vector(0 to 7) := (others => '0');
    variable r3169 : std_logic_vector(0 to 0) := (others => '0');
    variable r3167 : std_logic_vector(0 to 0) := (others => '0');
    variable r3165 : std_logic_vector(0 to 0) := (others => '0');
    variable r3163 : std_logic_vector(0 to 0) := (others => '0');
    variable r3161 : std_logic_vector(0 to 0) := (others => '0');
    variable r3159 : std_logic_vector(0 to 0) := (others => '0');
    variable r3157 : std_logic_vector(0 to 0) := (others => '0');
    variable r3155 : std_logic_vector(0 to 0) := (others => '0');
    variable r3153 : std_logic_vector(0 to 7) := (others => '0');
    variable r3151 : std_logic_vector(0 to 0) := (others => '0');
    variable r3149 : std_logic_vector(0 to 0) := (others => '0');
    variable r3147 : std_logic_vector(0 to 0) := (others => '0');
    variable r3145 : std_logic_vector(0 to 0) := (others => '0');
    variable r3143 : std_logic_vector(0 to 0) := (others => '0');
    variable r3141 : std_logic_vector(0 to 0) := (others => '0');
    variable r3139 : std_logic_vector(0 to 0) := (others => '0');
    variable r3137 : std_logic_vector(0 to 0) := (others => '0');
    variable r3135 : std_logic_vector(0 to 7) := (others => '0');
    variable r3133 : std_logic_vector(0 to 0) := (others => '0');
    variable r3131 : std_logic_vector(0 to 0) := (others => '0');
    variable r3129 : std_logic_vector(0 to 0) := (others => '0');
    variable r3127 : std_logic_vector(0 to 0) := (others => '0');
    variable r3125 : std_logic_vector(0 to 0) := (others => '0');
    variable r3123 : std_logic_vector(0 to 0) := (others => '0');
    variable r3121 : std_logic_vector(0 to 0) := (others => '0');
    variable r3119 : std_logic_vector(0 to 0) := (others => '0');
    variable r3117 : std_logic_vector(0 to 7) := (others => '0');
    variable r3115 : std_logic_vector(0 to 0) := (others => '0');
    variable r3113 : std_logic_vector(0 to 0) := (others => '0');
    variable r3111 : std_logic_vector(0 to 0) := (others => '0');
    variable r3109 : std_logic_vector(0 to 0) := (others => '0');
    variable r3107 : std_logic_vector(0 to 0) := (others => '0');
    variable r3105 : std_logic_vector(0 to 0) := (others => '0');
    variable r3103 : std_logic_vector(0 to 0) := (others => '0');
    variable r3101 : std_logic_vector(0 to 0) := (others => '0');
    variable r3099 : std_logic_vector(0 to 7) := (others => '0');
    variable r3097 : std_logic_vector(0 to 0) := (others => '0');
    variable r3095 : std_logic_vector(0 to 0) := (others => '0');
    variable r3093 : std_logic_vector(0 to 0) := (others => '0');
    variable r3091 : std_logic_vector(0 to 0) := (others => '0');
    variable r3089 : std_logic_vector(0 to 0) := (others => '0');
    variable r3087 : std_logic_vector(0 to 0) := (others => '0');
    variable r3085 : std_logic_vector(0 to 0) := (others => '0');
    variable r3083 : std_logic_vector(0 to 0) := (others => '0');
    variable r3081 : std_logic_vector(0 to 7) := (others => '0');
    variable r3079 : std_logic_vector(0 to 0) := (others => '0');
    variable r3077 : std_logic_vector(0 to 0) := (others => '0');
    variable r3075 : std_logic_vector(0 to 0) := (others => '0');
    variable r3073 : std_logic_vector(0 to 0) := (others => '0');
    variable r3071 : std_logic_vector(0 to 0) := (others => '0');
    variable r3069 : std_logic_vector(0 to 0) := (others => '0');
    variable r3067 : std_logic_vector(0 to 0) := (others => '0');
    variable r3065 : std_logic_vector(0 to 0) := (others => '0');
    variable r3063 : std_logic_vector(0 to 7) := (others => '0');
    variable r3061 : std_logic_vector(0 to 0) := (others => '0');
    variable r3059 : std_logic_vector(0 to 0) := (others => '0');
    variable r3057 : std_logic_vector(0 to 0) := (others => '0');
    variable r3055 : std_logic_vector(0 to 0) := (others => '0');
    variable r3053 : std_logic_vector(0 to 0) := (others => '0');
    variable r3051 : std_logic_vector(0 to 0) := (others => '0');
    variable r3049 : std_logic_vector(0 to 0) := (others => '0');
    variable r3047 : std_logic_vector(0 to 0) := (others => '0');
    variable r3045 : std_logic_vector(0 to 7) := (others => '0');
    variable r3043 : std_logic_vector(0 to 0) := (others => '0');
    variable r3041 : std_logic_vector(0 to 0) := (others => '0');
    variable r3039 : std_logic_vector(0 to 0) := (others => '0');
    variable r3037 : std_logic_vector(0 to 0) := (others => '0');
    variable r3035 : std_logic_vector(0 to 0) := (others => '0');
    variable r3033 : std_logic_vector(0 to 0) := (others => '0');
    variable r3031 : std_logic_vector(0 to 0) := (others => '0');
    variable r3029 : std_logic_vector(0 to 0) := (others => '0');
    variable r3027 : std_logic_vector(0 to 7) := (others => '0');
    variable r3025 : std_logic_vector(0 to 0) := (others => '0');
    variable r3023 : std_logic_vector(0 to 0) := (others => '0');
    variable r3021 : std_logic_vector(0 to 0) := (others => '0');
    variable r3019 : std_logic_vector(0 to 0) := (others => '0');
    variable r3017 : std_logic_vector(0 to 0) := (others => '0');
    variable r3015 : std_logic_vector(0 to 0) := (others => '0');
    variable r3013 : std_logic_vector(0 to 0) := (others => '0');
    variable r3011 : std_logic_vector(0 to 0) := (others => '0');
    variable r3009 : std_logic_vector(0 to 7) := (others => '0');
    variable r3007 : std_logic_vector(0 to 0) := (others => '0');
    variable r3005 : std_logic_vector(0 to 0) := (others => '0');
    variable r3003 : std_logic_vector(0 to 0) := (others => '0');
    variable r3001 : std_logic_vector(0 to 0) := (others => '0');
    variable r2999 : std_logic_vector(0 to 0) := (others => '0');
    variable r2997 : std_logic_vector(0 to 0) := (others => '0');
    variable r2995 : std_logic_vector(0 to 0) := (others => '0');
    variable r2993 : std_logic_vector(0 to 0) := (others => '0');
    variable r2991 : std_logic_vector(0 to 7) := (others => '0');
    variable r2989 : std_logic_vector(0 to 0) := (others => '0');
    variable r2987 : std_logic_vector(0 to 0) := (others => '0');
    variable r2985 : std_logic_vector(0 to 0) := (others => '0');
    variable r2983 : std_logic_vector(0 to 0) := (others => '0');
    variable r2981 : std_logic_vector(0 to 0) := (others => '0');
    variable r2979 : std_logic_vector(0 to 0) := (others => '0');
    variable r2977 : std_logic_vector(0 to 0) := (others => '0');
    variable r2975 : std_logic_vector(0 to 0) := (others => '0');
    variable r2973 : std_logic_vector(0 to 7) := (others => '0');
    variable r2971 : std_logic_vector(0 to 0) := (others => '0');
    variable r2969 : std_logic_vector(0 to 0) := (others => '0');
    variable r2967 : std_logic_vector(0 to 0) := (others => '0');
    variable r2965 : std_logic_vector(0 to 0) := (others => '0');
    variable r2963 : std_logic_vector(0 to 0) := (others => '0');
    variable r2961 : std_logic_vector(0 to 0) := (others => '0');
    variable r2959 : std_logic_vector(0 to 0) := (others => '0');
    variable r2957 : std_logic_vector(0 to 0) := (others => '0');
    variable r2955 : std_logic_vector(0 to 7) := (others => '0');
    variable r2953 : std_logic_vector(0 to 0) := (others => '0');
    variable r2951 : std_logic_vector(0 to 0) := (others => '0');
    variable r2949 : std_logic_vector(0 to 0) := (others => '0');
    variable r2947 : std_logic_vector(0 to 0) := (others => '0');
    variable r2945 : std_logic_vector(0 to 0) := (others => '0');
    variable r2943 : std_logic_vector(0 to 0) := (others => '0');
    variable r2941 : std_logic_vector(0 to 0) := (others => '0');
    variable r2939 : std_logic_vector(0 to 0) := (others => '0');
    variable EMPTY : std_logic_vector(0 to -1) := (others => '0');
  begin
    r2939 := "1";
    r2941 := "0";
    r2943 := "0";
    r2945 := "0";
    r2947 := "0";
    r2949 := "0";
    r2951 := "0";
    r2953 := "0";
    r2955 := (r2939 & r2941 & r2943 & r2945 & r2947 & r2949 & r2951 & r2953);
    r2957 := "0";
    r2959 := "1";
    r2961 := "0";
    r2963 := "0";
    r2965 := "0";
    r2967 := "0";
    r2969 := "0";
    r2971 := "0";
    r2973 := (r2957 & r2959 & r2961 & r2963 & r2965 & r2967 & r2969 & r2971);
    r2975 := "1";
    r2977 := "1";
    r2979 := "0";
    r2981 := "0";
    r2983 := "0";
    r2985 := "0";
    r2987 := "0";
    r2989 := "0";
    r2991 := (r2975 & r2977 & r2979 & r2981 & r2983 & r2985 & r2987 & r2989);
    r2993 := "0";
    r2995 := "0";
    r2997 := "1";
    r2999 := "0";
    r3001 := "0";
    r3003 := "0";
    r3005 := "0";
    r3007 := "0";
    r3009 := (r2993 & r2995 & r2997 & r2999 & r3001 & r3003 & r3005 & r3007);
    r3011 := "1";
    r3013 := "0";
    r3015 := "1";
    r3017 := "0";
    r3019 := "0";
    r3021 := "0";
    r3023 := "0";
    r3025 := "0";
    r3027 := (r3011 & r3013 & r3015 & r3017 & r3019 & r3021 & r3023 & r3025);
    r3029 := "0";
    r3031 := "1";
    r3033 := "1";
    r3035 := "0";
    r3037 := "0";
    r3039 := "0";
    r3041 := "0";
    r3043 := "0";
    r3045 := (r3029 & r3031 & r3033 & r3035 & r3037 & r3039 & r3041 & r3043);
    r3047 := "1";
    r3049 := "1";
    r3051 := "1";
    r3053 := "0";
    r3055 := "0";
    r3057 := "0";
    r3059 := "0";
    r3061 := "0";
    r3063 := (r3047 & r3049 & r3051 & r3053 & r3055 & r3057 & r3059 & r3061);
    r3065 := "0";
    r3067 := "0";
    r3069 := "0";
    r3071 := "1";
    r3073 := "0";
    r3075 := "0";
    r3077 := "0";
    r3079 := "0";
    r3081 := (r3065 & r3067 & r3069 & r3071 & r3073 & r3075 & r3077 & r3079);
    r3083 := "1";
    r3085 := "0";
    r3087 := "0";
    r3089 := "1";
    r3091 := "0";
    r3093 := "0";
    r3095 := "0";
    r3097 := "0";
    r3099 := (r3083 & r3085 & r3087 & r3089 & r3091 & r3093 & r3095 & r3097);
    r3101 := "0";
    r3103 := "1";
    r3105 := "0";
    r3107 := "1";
    r3109 := "0";
    r3111 := "0";
    r3113 := "0";
    r3115 := "0";
    r3117 := (r3101 & r3103 & r3105 & r3107 & r3109 & r3111 & r3113 & r3115);
    r3119 := "1";
    r3121 := "1";
    r3123 := "0";
    r3125 := "1";
    r3127 := "0";
    r3129 := "0";
    r3131 := "0";
    r3133 := "0";
    r3135 := (r3119 & r3121 & r3123 & r3125 & r3127 & r3129 & r3131 & r3133);
    r3137 := "0";
    r3139 := "0";
    r3141 := "1";
    r3143 := "1";
    r3145 := "0";
    r3147 := "0";
    r3149 := "0";
    r3151 := "0";
    r3153 := (r3137 & r3139 & r3141 & r3143 & r3145 & r3147 & r3149 & r3151);
    r3155 := "1";
    r3157 := "0";
    r3159 := "1";
    r3161 := "1";
    r3163 := "0";
    r3165 := "0";
    r3167 := "0";
    r3169 := "0";
    r3171 := (r3155 & r3157 & r3159 & r3161 & r3163 & r3165 & r3167 & r3169);
    r3173 := "0";
    r3175 := "1";
    r3177 := "1";
    r3179 := "1";
    r3181 := "0";
    r3183 := "0";
    r3185 := "0";
    r3187 := "0";
    r3189 := (r3173 & r3175 & r3177 & r3179 & r3181 & r3183 & r3185 & r3187);
    r3191 := "1";
    r3193 := "1";
    r3195 := "1";
    r3197 := "1";
    r3199 := "0";
    r3201 := "0";
    r3203 := "0";
    r3205 := "0";
    r3207 := (r3191 & r3193 & r3195 & r3197 & r3199 & r3201 & r3203 & r3205);
    r3209 := "0";
    r3211 := "0";
    r3213 := "0";
    r3215 := "0";
    r3217 := "1";
    r3219 := "0";
    r3221 := "0";
    r3223 := "0";
    r3225 := (r3209 & r3211 & r3213 & r3215 & r3217 & r3219 & r3221 & r3223);
    r3226 := (r2955 & r2973 & r2991 & r3009 & r3027 & r3045 & r3063 & r3081 & r3099 & r3117 & r3135 & r3153 & r3171 & r3189 & r3207 & r3225);
    return r3226;
  end rewire_key1_2935;
  function rewire_buildSalsa256_1178(r1179 : std_logic_vector ; r1180 : std_logic_vector ; r1181 : std_logic_vector ; r1182 : std_logic_vector) return std_logic_vector
  is
    variable r2934 : std_logic_vector(0 to 511) := (others => '0');
    variable r2933 : std_logic_vector(0 to 511) := (others => '0');
    variable r1656 : std_logic_vector(0 to 511) := (others => '0');
    variable r1655 : std_logic_vector(0 to 511) := (others => '0');
    variable b1653 : boolean := false;
    variable b1652 : boolean := false;
    variable b1651 : boolean := false;
    variable b1650 : boolean := false;
    variable b1649 : boolean := false;
    variable b1648 : boolean := false;
    variable r1647 : std_logic_vector(0 to 7) := (others => '0');
    variable r1646 : std_logic_vector(0 to 7) := (others => '0');
    variable r1645 : std_logic_vector(0 to 7) := (others => '0');
    variable r1644 : std_logic_vector(0 to 7) := (others => '0');
    variable b1643 : boolean := false;
    variable b1642 : boolean := false;
    variable b1641 : boolean := false;
    variable b1640 : boolean := false;
    variable b1639 : boolean := false;
    variable b1638 : boolean := false;
    variable r1637 : std_logic_vector(0 to 7) := (others => '0');
    variable r1636 : std_logic_vector(0 to 7) := (others => '0');
    variable r1635 : std_logic_vector(0 to 7) := (others => '0');
    variable r1634 : std_logic_vector(0 to 7) := (others => '0');
    variable b1633 : boolean := false;
    variable b1632 : boolean := false;
    variable b1631 : boolean := false;
    variable b1630 : boolean := false;
    variable b1629 : boolean := false;
    variable b1628 : boolean := false;
    variable r1627 : std_logic_vector(0 to 7) := (others => '0');
    variable r1626 : std_logic_vector(0 to 7) := (others => '0');
    variable r1625 : std_logic_vector(0 to 7) := (others => '0');
    variable r1624 : std_logic_vector(0 to 7) := (others => '0');
    variable b1623 : boolean := false;
    variable b1622 : boolean := false;
    variable b1621 : boolean := false;
    variable b1620 : boolean := false;
    variable b1619 : boolean := false;
    variable b1618 : boolean := false;
    variable r1617 : std_logic_vector(0 to 7) := (others => '0');
    variable r1616 : std_logic_vector(0 to 7) := (others => '0');
    variable r1615 : std_logic_vector(0 to 7) := (others => '0');
    variable r1614 : std_logic_vector(0 to 7) := (others => '0');
    variable b1613 : boolean := false;
    variable r1612 : std_logic_vector(0 to 31) := (others => '0');
    variable r1611 : std_logic_vector(0 to 31) := (others => '0');
    variable r1610 : std_logic_vector(0 to 31) := (others => '0');
    variable r1609 : std_logic_vector(0 to 31) := (others => '0');
    variable b1608 : boolean := false;
    variable r1607 : std_logic_vector(0 to 511) := (others => '0');
    variable r1606 : std_logic_vector(0 to 127) := (others => '0');
    variable r1605 : std_logic_vector(0 to 31) := (others => '0');
    variable r1530 : std_logic_vector(0 to 31) := (others => '0');
    variable r1528 : std_logic_vector(0 to 31) := (others => '0');
    variable r1453 : std_logic_vector(0 to 31) := (others => '0');
    variable r1451 : std_logic_vector(0 to 31) := (others => '0');
    variable r1376 : std_logic_vector(0 to 31) := (others => '0');
    variable r1374 : std_logic_vector(0 to 31) := (others => '0');
    variable r1299 : std_logic_vector(0 to 31) := (others => '0');
    variable b1296 : boolean := false;
    variable b1295 : boolean := false;
    variable b1294 : boolean := false;
    variable b1293 : boolean := false;
    variable b1292 : boolean := false;
    variable b1291 : boolean := false;
    variable b1290 : boolean := false;
    variable b1289 : boolean := false;
    variable b1288 : boolean := false;
    variable b1287 : boolean := false;
    variable r1286 : std_logic_vector(0 to 7) := (others => '0');
    variable r1285 : std_logic_vector(0 to 7) := (others => '0');
    variable r1284 : std_logic_vector(0 to 7) := (others => '0');
    variable r1283 : std_logic_vector(0 to 7) := (others => '0');
    variable r1282 : std_logic_vector(0 to 7) := (others => '0');
    variable r1281 : std_logic_vector(0 to 7) := (others => '0');
    variable r1280 : std_logic_vector(0 to 7) := (others => '0');
    variable r1279 : std_logic_vector(0 to 7) := (others => '0');
    variable b1278 : boolean := false;
    variable b1277 : boolean := false;
    variable b1276 : boolean := false;
    variable b1275 : boolean := false;
    variable b1274 : boolean := false;
    variable b1273 : boolean := false;
    variable b1272 : boolean := false;
    variable b1271 : boolean := false;
    variable b1270 : boolean := false;
    variable b1269 : boolean := false;
    variable r1268 : std_logic_vector(0 to 7) := (others => '0');
    variable r1267 : std_logic_vector(0 to 7) := (others => '0');
    variable r1266 : std_logic_vector(0 to 7) := (others => '0');
    variable r1265 : std_logic_vector(0 to 7) := (others => '0');
    variable r1264 : std_logic_vector(0 to 7) := (others => '0');
    variable r1263 : std_logic_vector(0 to 7) := (others => '0');
    variable r1262 : std_logic_vector(0 to 7) := (others => '0');
    variable r1261 : std_logic_vector(0 to 7) := (others => '0');
    variable b1260 : boolean := false;
    variable b1259 : boolean := false;
    variable b1258 : boolean := false;
    variable b1257 : boolean := false;
    variable b1256 : boolean := false;
    variable b1255 : boolean := false;
    variable b1254 : boolean := false;
    variable b1253 : boolean := false;
    variable b1252 : boolean := false;
    variable b1251 : boolean := false;
    variable b1250 : boolean := false;
    variable b1249 : boolean := false;
    variable b1248 : boolean := false;
    variable b1247 : boolean := false;
    variable b1246 : boolean := false;
    variable b1245 : boolean := false;
    variable b1244 : boolean := false;
    variable b1243 : boolean := false;
    variable r1242 : std_logic_vector(0 to 7) := (others => '0');
    variable r1241 : std_logic_vector(0 to 7) := (others => '0');
    variable r1240 : std_logic_vector(0 to 7) := (others => '0');
    variable r1239 : std_logic_vector(0 to 7) := (others => '0');
    variable r1238 : std_logic_vector(0 to 7) := (others => '0');
    variable r1237 : std_logic_vector(0 to 7) := (others => '0');
    variable r1236 : std_logic_vector(0 to 7) := (others => '0');
    variable r1235 : std_logic_vector(0 to 7) := (others => '0');
    variable r1234 : std_logic_vector(0 to 7) := (others => '0');
    variable r1233 : std_logic_vector(0 to 7) := (others => '0');
    variable r1232 : std_logic_vector(0 to 7) := (others => '0');
    variable r1231 : std_logic_vector(0 to 7) := (others => '0');
    variable r1230 : std_logic_vector(0 to 7) := (others => '0');
    variable r1229 : std_logic_vector(0 to 7) := (others => '0');
    variable r1228 : std_logic_vector(0 to 7) := (others => '0');
    variable r1227 : std_logic_vector(0 to 7) := (others => '0');
    variable b1226 : boolean := false;
    variable b1225 : boolean := false;
    variable b1224 : boolean := false;
    variable b1223 : boolean := false;
    variable b1222 : boolean := false;
    variable b1221 : boolean := false;
    variable b1220 : boolean := false;
    variable b1219 : boolean := false;
    variable b1218 : boolean := false;
    variable b1217 : boolean := false;
    variable b1216 : boolean := false;
    variable b1215 : boolean := false;
    variable b1214 : boolean := false;
    variable b1213 : boolean := false;
    variable b1212 : boolean := false;
    variable b1211 : boolean := false;
    variable b1210 : boolean := false;
    variable b1209 : boolean := false;
    variable r1208 : std_logic_vector(0 to 7) := (others => '0');
    variable r1207 : std_logic_vector(0 to 7) := (others => '0');
    variable r1206 : std_logic_vector(0 to 7) := (others => '0');
    variable r1205 : std_logic_vector(0 to 7) := (others => '0');
    variable r1204 : std_logic_vector(0 to 7) := (others => '0');
    variable r1203 : std_logic_vector(0 to 7) := (others => '0');
    variable r1202 : std_logic_vector(0 to 7) := (others => '0');
    variable r1201 : std_logic_vector(0 to 7) := (others => '0');
    variable r1200 : std_logic_vector(0 to 7) := (others => '0');
    variable r1199 : std_logic_vector(0 to 7) := (others => '0');
    variable r1198 : std_logic_vector(0 to 7) := (others => '0');
    variable r1197 : std_logic_vector(0 to 7) := (others => '0');
    variable r1196 : std_logic_vector(0 to 7) := (others => '0');
    variable r1195 : std_logic_vector(0 to 7) := (others => '0');
    variable r1194 : std_logic_vector(0 to 7) := (others => '0');
    variable r1193 : std_logic_vector(0 to 7) := (others => '0');
    variable b1192 : boolean := false;
    variable r1191 : std_logic_vector(0 to 63) := (others => '0');
    variable r1190 : std_logic_vector(0 to 63) := (others => '0');
    variable r1189 : std_logic_vector(0 to 127) := (others => '0');
    variable r1188 : std_logic_vector(0 to 127) := (others => '0');
    variable b1187 : boolean := false;
    variable r1186 : std_logic_vector(0 to 511) := (others => '0');
    variable r1185 : std_logic_vector(0 to 383) := (others => '0');
    variable EMPTY : std_logic_vector(0 to -1) := (others => '0');
  begin
    b1187 := true;
    r1188 := r1185(0 to 127);
    r1189 := r1185(128 to 255);
    r1190 := r1185(256 to 319);
    r1191 := r1185(320 to 383);
    b1192 := true;
    r1193 := r1188(0 to 7);
    r1194 := r1188(8 to 15);
    r1195 := r1188(16 to 23);
    r1196 := r1188(24 to 31);
    r1197 := r1188(32 to 39);
    r1198 := r1188(40 to 47);
    r1199 := r1188(48 to 55);
    r1200 := r1188(56 to 63);
    r1201 := r1188(64 to 71);
    r1202 := r1188(72 to 79);
    r1203 := r1188(80 to 87);
    r1204 := r1188(88 to 95);
    r1205 := r1188(96 to 103);
    r1206 := r1188(104 to 111);
    r1207 := r1188(112 to 119);
    r1208 := r1188(120 to 127);
    b1209 := true;
    b1210 := true;
    b1211 := true;
    b1212 := true;
    b1213 := true;
    b1214 := true;
    b1215 := true;
    b1216 := true;
    b1217 := true;
    b1218 := true;
    b1219 := true;
    b1220 := true;
    b1221 := true;
    b1222 := true;
    b1223 := true;
    b1224 := true;
    b1225 := (b1209 AND (b1210 AND (b1211 AND (b1212 AND (b1213 AND (b1214 AND (b1215 AND (b1216 AND (b1217 AND (b1218 AND (b1219 AND (b1220 AND (b1221 AND (b1222 AND (b1223 AND b1224)))))))))))))));
    b1226 := true;
    r1227 := r1189(0 to 7);
    r1228 := r1189(8 to 15);
    r1229 := r1189(16 to 23);
    r1230 := r1189(24 to 31);
    r1231 := r1189(32 to 39);
    r1232 := r1189(40 to 47);
    r1233 := r1189(48 to 55);
    r1234 := r1189(56 to 63);
    r1235 := r1189(64 to 71);
    r1236 := r1189(72 to 79);
    r1237 := r1189(80 to 87);
    r1238 := r1189(88 to 95);
    r1239 := r1189(96 to 103);
    r1240 := r1189(104 to 111);
    r1241 := r1189(112 to 119);
    r1242 := r1189(120 to 127);
    b1243 := true;
    b1244 := true;
    b1245 := true;
    b1246 := true;
    b1247 := true;
    b1248 := true;
    b1249 := true;
    b1250 := true;
    b1251 := true;
    b1252 := true;
    b1253 := true;
    b1254 := true;
    b1255 := true;
    b1256 := true;
    b1257 := true;
    b1258 := true;
    b1259 := (b1243 AND (b1244 AND (b1245 AND (b1246 AND (b1247 AND (b1248 AND (b1249 AND (b1250 AND (b1251 AND (b1252 AND (b1253 AND (b1254 AND (b1255 AND (b1256 AND (b1257 AND b1258)))))))))))))));
    b1260 := true;
    r1261 := r1190(0 to 7);
    r1262 := r1190(8 to 15);
    r1263 := r1190(16 to 23);
    r1264 := r1190(24 to 31);
    r1265 := r1190(32 to 39);
    r1266 := r1190(40 to 47);
    r1267 := r1190(48 to 55);
    r1268 := r1190(56 to 63);
    b1269 := true;
    b1270 := true;
    b1271 := true;
    b1272 := true;
    b1273 := true;
    b1274 := true;
    b1275 := true;
    b1276 := true;
    b1277 := (b1269 AND (b1270 AND (b1271 AND (b1272 AND (b1273 AND (b1274 AND (b1275 AND b1276)))))));
    b1278 := true;
    r1279 := r1191(0 to 7);
    r1280 := r1191(8 to 15);
    r1281 := r1191(16 to 23);
    r1282 := r1191(24 to 31);
    r1283 := r1191(32 to 39);
    r1284 := r1191(40 to 47);
    r1285 := r1191(48 to 55);
    r1286 := r1191(56 to 63);
    b1287 := true;
    b1288 := true;
    b1289 := true;
    b1290 := true;
    b1291 := true;
    b1292 := true;
    b1293 := true;
    b1294 := true;
    b1295 := (b1287 AND (b1288 AND (b1289 AND (b1290 AND (b1291 AND (b1292 AND (b1293 AND b1294)))))));
    b1296 := (b1225 AND (b1259 AND (b1277 AND b1295)));
    if b1296 then
      b1608 := true;
      r1609 := r1606(0 to 31);
      r1610 := r1606(32 to 63);
      r1611 := r1606(64 to 95);
      r1612 := r1606(96 to 127);
      b1613 := true;
      r1614 := r1609(0 to 7);
      r1615 := r1609(8 to 15);
      r1616 := r1609(16 to 23);
      r1617 := r1609(24 to 31);
      b1618 := true;
      b1619 := true;
      b1620 := true;
      b1621 := true;
      b1622 := (b1618 AND (b1619 AND (b1620 AND b1621)));
      b1623 := true;
      r1624 := r1610(0 to 7);
      r1625 := r1610(8 to 15);
      r1626 := r1610(16 to 23);
      r1627 := r1610(24 to 31);
      b1628 := true;
      b1629 := true;
      b1630 := true;
      b1631 := true;
      b1632 := (b1628 AND (b1629 AND (b1630 AND b1631)));
      b1633 := true;
      r1634 := r1611(0 to 7);
      r1635 := r1611(8 to 15);
      r1636 := r1611(16 to 23);
      r1637 := r1611(24 to 31);
      b1638 := true;
      b1639 := true;
      b1640 := true;
      b1641 := true;
      b1642 := (b1638 AND (b1639 AND (b1640 AND b1641)));
      b1643 := true;
      r1644 := r1612(0 to 7);
      r1645 := r1612(8 to 15);
      r1646 := r1612(16 to 23);
      r1647 := r1612(24 to 31);
      b1648 := true;
      b1649 := true;
      b1650 := true;
      b1651 := true;
      b1652 := (b1648 AND (b1649 AND (b1650 AND b1651)));
      b1653 := (b1622 AND (b1632 AND (b1642 AND b1652)));
      if b1653 then
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        r2933 := (r1614 & r1615 & r1616 & r1617 & r1193 & r1194 & r1195 & r1196 & r1197 & r1198 & r1199 & r1200 & r1201 & r1202 & r1203 & r1204 & r1205 & r1206 & r1207 & r1208 & r1624 & r1625 & r1626 & r1627 & r1261 & r1262 & r1263 & r1264 & r1265 & r1266 & r1267 & r1268 & r1279 & r1280 & r1281 & r1282 & r1283 & r1284 & r1285 & r1286 & r1634 & r1635 & r1636 & r1637 & r1227 & r1228 & r1229 & r1230 & r1231 & r1232 & r1233 & r1234 & r1235 & r1236 & r1237 & r1238 & r1239 & r1240 & r1241 & r1242 & r1644 & r1645 & r1646 & r1647);
        r2934 := rewire_salsaHash_1654(r2933);
        r1607 := r2934;
      end if;
      r1186 := r1607;
    end if;
    return r1186;
  end rewire_buildSalsa256_1178;
  function rewire_salsaHash_1654(r1655 : std_logic_vector) return std_logic_vector
  is
    variable r2931 : std_logic_vector(0 to 511) := (others => '0');
    variable r2930 : std_logic_vector(0 to 511) := (others => '0');
    variable r2929 : std_logic_vector(0 to 511) := (others => '0');
    variable r2600 : std_logic_vector(0 to 511) := (others => '0');
    variable r2599 : std_logic_vector(0 to 511) := (others => '0');
    variable r1976 : std_logic_vector(0 to 511) := (others => '0');
    variable r1975 : std_logic_vector(0 to 511) := (others => '0');
    variable r1659 : std_logic_vector(0 to 511) := (others => '0');
    variable r1658 : std_logic_vector(0 to 511) := (others => '0');
  begin
    null;
    r2929 := rewire_impwords_2598(r1655);
    r2930 := rewire_salsaHashp_1974(r2929);
    r2931 := rewire_expwords_1657(r2930);
    return r2931;
  end rewire_salsaHash_1654;
  function rewire_impwords_2598(r2599 : std_logic_vector) return std_logic_vector
  is
    variable r2928 : std_logic_vector(0 to 511) := (others => '0');
    variable r2926 : std_logic_vector(0 to 31) := (others => '0');
    variable r2925 : std_logic_vector(0 to 31) := (others => '0');
    variable r2923 : std_logic_vector(0 to 31) := (others => '0');
    variable r2922 : std_logic_vector(0 to 31) := (others => '0');
    variable r2920 : std_logic_vector(0 to 31) := (others => '0');
    variable r2919 : std_logic_vector(0 to 31) := (others => '0');
    variable r2917 : std_logic_vector(0 to 31) := (others => '0');
    variable r2916 : std_logic_vector(0 to 31) := (others => '0');
    variable r2914 : std_logic_vector(0 to 31) := (others => '0');
    variable r2913 : std_logic_vector(0 to 31) := (others => '0');
    variable r2911 : std_logic_vector(0 to 31) := (others => '0');
    variable r2910 : std_logic_vector(0 to 31) := (others => '0');
    variable r2908 : std_logic_vector(0 to 31) := (others => '0');
    variable r2907 : std_logic_vector(0 to 31) := (others => '0');
    variable r2905 : std_logic_vector(0 to 31) := (others => '0');
    variable r2904 : std_logic_vector(0 to 31) := (others => '0');
    variable r2902 : std_logic_vector(0 to 31) := (others => '0');
    variable r2901 : std_logic_vector(0 to 31) := (others => '0');
    variable r2899 : std_logic_vector(0 to 31) := (others => '0');
    variable r2898 : std_logic_vector(0 to 31) := (others => '0');
    variable r2896 : std_logic_vector(0 to 31) := (others => '0');
    variable r2895 : std_logic_vector(0 to 31) := (others => '0');
    variable r2893 : std_logic_vector(0 to 31) := (others => '0');
    variable r2892 : std_logic_vector(0 to 31) := (others => '0');
    variable r2890 : std_logic_vector(0 to 31) := (others => '0');
    variable r2889 : std_logic_vector(0 to 31) := (others => '0');
    variable r2887 : std_logic_vector(0 to 31) := (others => '0');
    variable r2886 : std_logic_vector(0 to 31) := (others => '0');
    variable r2884 : std_logic_vector(0 to 31) := (others => '0');
    variable r2883 : std_logic_vector(0 to 31) := (others => '0');
    variable r2881 : std_logic_vector(0 to 31) := (others => '0');
    variable r2880 : std_logic_vector(0 to 31) := (others => '0');
    variable EMPTY : std_logic_vector(0 to -1) := (others => '0');
    variable r2734 : std_logic_vector(0 to 31) := (others => '0');
    variable r2733 : std_logic_vector(0 to 31) := (others => '0');
    variable b2731 : boolean := false;
    variable b2730 : boolean := false;
    variable b2729 : boolean := false;
    variable b2728 : boolean := false;
    variable b2727 : boolean := false;
    variable b2726 : boolean := false;
    variable b2725 : boolean := false;
    variable b2724 : boolean := false;
    variable b2723 : boolean := false;
    variable b2722 : boolean := false;
    variable b2721 : boolean := false;
    variable b2720 : boolean := false;
    variable b2719 : boolean := false;
    variable b2718 : boolean := false;
    variable b2717 : boolean := false;
    variable b2716 : boolean := false;
    variable b2715 : boolean := false;
    variable b2714 : boolean := false;
    variable b2713 : boolean := false;
    variable b2712 : boolean := false;
    variable b2711 : boolean := false;
    variable b2710 : boolean := false;
    variable b2709 : boolean := false;
    variable b2708 : boolean := false;
    variable b2707 : boolean := false;
    variable b2706 : boolean := false;
    variable b2705 : boolean := false;
    variable b2704 : boolean := false;
    variable b2703 : boolean := false;
    variable b2702 : boolean := false;
    variable b2701 : boolean := false;
    variable b2700 : boolean := false;
    variable b2699 : boolean := false;
    variable b2698 : boolean := false;
    variable b2697 : boolean := false;
    variable b2696 : boolean := false;
    variable b2695 : boolean := false;
    variable b2694 : boolean := false;
    variable b2693 : boolean := false;
    variable b2692 : boolean := false;
    variable b2691 : boolean := false;
    variable b2690 : boolean := false;
    variable b2689 : boolean := false;
    variable b2688 : boolean := false;
    variable b2687 : boolean := false;
    variable b2686 : boolean := false;
    variable b2685 : boolean := false;
    variable b2684 : boolean := false;
    variable b2683 : boolean := false;
    variable b2682 : boolean := false;
    variable b2681 : boolean := false;
    variable b2680 : boolean := false;
    variable b2679 : boolean := false;
    variable b2678 : boolean := false;
    variable b2677 : boolean := false;
    variable b2676 : boolean := false;
    variable b2675 : boolean := false;
    variable b2674 : boolean := false;
    variable b2673 : boolean := false;
    variable b2672 : boolean := false;
    variable b2671 : boolean := false;
    variable b2670 : boolean := false;
    variable b2669 : boolean := false;
    variable b2668 : boolean := false;
    variable b2667 : boolean := false;
    variable r2666 : std_logic_vector(0 to 7) := (others => '0');
    variable r2665 : std_logic_vector(0 to 7) := (others => '0');
    variable r2664 : std_logic_vector(0 to 7) := (others => '0');
    variable r2663 : std_logic_vector(0 to 7) := (others => '0');
    variable r2662 : std_logic_vector(0 to 7) := (others => '0');
    variable r2661 : std_logic_vector(0 to 7) := (others => '0');
    variable r2660 : std_logic_vector(0 to 7) := (others => '0');
    variable r2659 : std_logic_vector(0 to 7) := (others => '0');
    variable r2658 : std_logic_vector(0 to 7) := (others => '0');
    variable r2657 : std_logic_vector(0 to 7) := (others => '0');
    variable r2656 : std_logic_vector(0 to 7) := (others => '0');
    variable r2655 : std_logic_vector(0 to 7) := (others => '0');
    variable r2654 : std_logic_vector(0 to 7) := (others => '0');
    variable r2653 : std_logic_vector(0 to 7) := (others => '0');
    variable r2652 : std_logic_vector(0 to 7) := (others => '0');
    variable r2651 : std_logic_vector(0 to 7) := (others => '0');
    variable r2650 : std_logic_vector(0 to 7) := (others => '0');
    variable r2649 : std_logic_vector(0 to 7) := (others => '0');
    variable r2648 : std_logic_vector(0 to 7) := (others => '0');
    variable r2647 : std_logic_vector(0 to 7) := (others => '0');
    variable r2646 : std_logic_vector(0 to 7) := (others => '0');
    variable r2645 : std_logic_vector(0 to 7) := (others => '0');
    variable r2644 : std_logic_vector(0 to 7) := (others => '0');
    variable r2643 : std_logic_vector(0 to 7) := (others => '0');
    variable r2642 : std_logic_vector(0 to 7) := (others => '0');
    variable r2641 : std_logic_vector(0 to 7) := (others => '0');
    variable r2640 : std_logic_vector(0 to 7) := (others => '0');
    variable r2639 : std_logic_vector(0 to 7) := (others => '0');
    variable r2638 : std_logic_vector(0 to 7) := (others => '0');
    variable r2637 : std_logic_vector(0 to 7) := (others => '0');
    variable r2636 : std_logic_vector(0 to 7) := (others => '0');
    variable r2635 : std_logic_vector(0 to 7) := (others => '0');
    variable r2634 : std_logic_vector(0 to 7) := (others => '0');
    variable r2633 : std_logic_vector(0 to 7) := (others => '0');
    variable r2632 : std_logic_vector(0 to 7) := (others => '0');
    variable r2631 : std_logic_vector(0 to 7) := (others => '0');
    variable r2630 : std_logic_vector(0 to 7) := (others => '0');
    variable r2629 : std_logic_vector(0 to 7) := (others => '0');
    variable r2628 : std_logic_vector(0 to 7) := (others => '0');
    variable r2627 : std_logic_vector(0 to 7) := (others => '0');
    variable r2626 : std_logic_vector(0 to 7) := (others => '0');
    variable r2625 : std_logic_vector(0 to 7) := (others => '0');
    variable r2624 : std_logic_vector(0 to 7) := (others => '0');
    variable r2623 : std_logic_vector(0 to 7) := (others => '0');
    variable r2622 : std_logic_vector(0 to 7) := (others => '0');
    variable r2621 : std_logic_vector(0 to 7) := (others => '0');
    variable r2620 : std_logic_vector(0 to 7) := (others => '0');
    variable r2619 : std_logic_vector(0 to 7) := (others => '0');
    variable r2618 : std_logic_vector(0 to 7) := (others => '0');
    variable r2617 : std_logic_vector(0 to 7) := (others => '0');
    variable r2616 : std_logic_vector(0 to 7) := (others => '0');
    variable r2615 : std_logic_vector(0 to 7) := (others => '0');
    variable r2614 : std_logic_vector(0 to 7) := (others => '0');
    variable r2613 : std_logic_vector(0 to 7) := (others => '0');
    variable r2612 : std_logic_vector(0 to 7) := (others => '0');
    variable r2611 : std_logic_vector(0 to 7) := (others => '0');
    variable r2610 : std_logic_vector(0 to 7) := (others => '0');
    variable r2609 : std_logic_vector(0 to 7) := (others => '0');
    variable r2608 : std_logic_vector(0 to 7) := (others => '0');
    variable r2607 : std_logic_vector(0 to 7) := (others => '0');
    variable r2606 : std_logic_vector(0 to 7) := (others => '0');
    variable r2605 : std_logic_vector(0 to 7) := (others => '0');
    variable r2604 : std_logic_vector(0 to 7) := (others => '0');
    variable r2603 : std_logic_vector(0 to 7) := (others => '0');
    variable b2602 : boolean := false;
    variable r2601 : std_logic_vector(0 to 511) := (others => '0');
  begin
    b2602 := true;
    r2603 := r2599(0 to 7);
    r2604 := r2599(8 to 15);
    r2605 := r2599(16 to 23);
    r2606 := r2599(24 to 31);
    r2607 := r2599(32 to 39);
    r2608 := r2599(40 to 47);
    r2609 := r2599(48 to 55);
    r2610 := r2599(56 to 63);
    r2611 := r2599(64 to 71);
    r2612 := r2599(72 to 79);
    r2613 := r2599(80 to 87);
    r2614 := r2599(88 to 95);
    r2615 := r2599(96 to 103);
    r2616 := r2599(104 to 111);
    r2617 := r2599(112 to 119);
    r2618 := r2599(120 to 127);
    r2619 := r2599(128 to 135);
    r2620 := r2599(136 to 143);
    r2621 := r2599(144 to 151);
    r2622 := r2599(152 to 159);
    r2623 := r2599(160 to 167);
    r2624 := r2599(168 to 175);
    r2625 := r2599(176 to 183);
    r2626 := r2599(184 to 191);
    r2627 := r2599(192 to 199);
    r2628 := r2599(200 to 207);
    r2629 := r2599(208 to 215);
    r2630 := r2599(216 to 223);
    r2631 := r2599(224 to 231);
    r2632 := r2599(232 to 239);
    r2633 := r2599(240 to 247);
    r2634 := r2599(248 to 255);
    r2635 := r2599(256 to 263);
    r2636 := r2599(264 to 271);
    r2637 := r2599(272 to 279);
    r2638 := r2599(280 to 287);
    r2639 := r2599(288 to 295);
    r2640 := r2599(296 to 303);
    r2641 := r2599(304 to 311);
    r2642 := r2599(312 to 319);
    r2643 := r2599(320 to 327);
    r2644 := r2599(328 to 335);
    r2645 := r2599(336 to 343);
    r2646 := r2599(344 to 351);
    r2647 := r2599(352 to 359);
    r2648 := r2599(360 to 367);
    r2649 := r2599(368 to 375);
    r2650 := r2599(376 to 383);
    r2651 := r2599(384 to 391);
    r2652 := r2599(392 to 399);
    r2653 := r2599(400 to 407);
    r2654 := r2599(408 to 415);
    r2655 := r2599(416 to 423);
    r2656 := r2599(424 to 431);
    r2657 := r2599(432 to 439);
    r2658 := r2599(440 to 447);
    r2659 := r2599(448 to 455);
    r2660 := r2599(456 to 463);
    r2661 := r2599(464 to 471);
    r2662 := r2599(472 to 479);
    r2663 := r2599(480 to 487);
    r2664 := r2599(488 to 495);
    r2665 := r2599(496 to 503);
    r2666 := r2599(504 to 511);
    b2667 := true;
    b2668 := true;
    b2669 := true;
    b2670 := true;
    b2671 := true;
    b2672 := true;
    b2673 := true;
    b2674 := true;
    b2675 := true;
    b2676 := true;
    b2677 := true;
    b2678 := true;
    b2679 := true;
    b2680 := true;
    b2681 := true;
    b2682 := true;
    b2683 := true;
    b2684 := true;
    b2685 := true;
    b2686 := true;
    b2687 := true;
    b2688 := true;
    b2689 := true;
    b2690 := true;
    b2691 := true;
    b2692 := true;
    b2693 := true;
    b2694 := true;
    b2695 := true;
    b2696 := true;
    b2697 := true;
    b2698 := true;
    b2699 := true;
    b2700 := true;
    b2701 := true;
    b2702 := true;
    b2703 := true;
    b2704 := true;
    b2705 := true;
    b2706 := true;
    b2707 := true;
    b2708 := true;
    b2709 := true;
    b2710 := true;
    b2711 := true;
    b2712 := true;
    b2713 := true;
    b2714 := true;
    b2715 := true;
    b2716 := true;
    b2717 := true;
    b2718 := true;
    b2719 := true;
    b2720 := true;
    b2721 := true;
    b2722 := true;
    b2723 := true;
    b2724 := true;
    b2725 := true;
    b2726 := true;
    b2727 := true;
    b2728 := true;
    b2729 := true;
    b2730 := true;
    b2731 := (b2667 AND (b2668 AND (b2669 AND (b2670 AND (b2671 AND (b2672 AND (b2673 AND (b2674 AND (b2675 AND (b2676 AND (b2677 AND (b2678 AND (b2679 AND (b2680 AND (b2681 AND (b2682 AND (b2683 AND (b2684 AND (b2685 AND (b2686 AND (b2687 AND (b2688 AND (b2689 AND (b2690 AND (b2691 AND (b2692 AND (b2693 AND (b2694 AND (b2695 AND (b2696 AND (b2697 AND (b2698 AND (b2699 AND (b2700 AND (b2701 AND (b2702 AND (b2703 AND (b2704 AND (b2705 AND (b2706 AND (b2707 AND (b2708 AND (b2709 AND (b2710 AND (b2711 AND (b2712 AND (b2713 AND (b2714 AND (b2715 AND (b2716 AND (b2717 AND (b2718 AND (b2719 AND (b2720 AND (b2721 AND (b2722 AND (b2723 AND (b2724 AND (b2725 AND (b2726 AND (b2727 AND (b2728 AND (b2729 AND b2730)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
    if b2731 then
      null;
      null;
      null;
      null;
      r2880 := (r2603 & r2604 & r2605 & r2606);
      r2881 := rewire_littleendian_2732(r2880);
      null;
      null;
      null;
      null;
      r2883 := (r2607 & r2608 & r2609 & r2610);
      r2884 := rewire_littleendian_2732(r2883);
      null;
      null;
      null;
      null;
      r2886 := (r2611 & r2612 & r2613 & r2614);
      r2887 := rewire_littleendian_2732(r2886);
      null;
      null;
      null;
      null;
      r2889 := (r2615 & r2616 & r2617 & r2618);
      r2890 := rewire_littleendian_2732(r2889);
      null;
      null;
      null;
      null;
      r2892 := (r2619 & r2620 & r2621 & r2622);
      r2893 := rewire_littleendian_2732(r2892);
      null;
      null;
      null;
      null;
      r2895 := (r2623 & r2624 & r2625 & r2626);
      r2896 := rewire_littleendian_2732(r2895);
      null;
      null;
      null;
      null;
      r2898 := (r2627 & r2628 & r2629 & r2630);
      r2899 := rewire_littleendian_2732(r2898);
      null;
      null;
      null;
      null;
      r2901 := (r2631 & r2632 & r2633 & r2634);
      r2902 := rewire_littleendian_2732(r2901);
      null;
      null;
      null;
      null;
      r2904 := (r2635 & r2636 & r2637 & r2638);
      r2905 := rewire_littleendian_2732(r2904);
      null;
      null;
      null;
      null;
      r2907 := (r2639 & r2640 & r2641 & r2642);
      r2908 := rewire_littleendian_2732(r2907);
      null;
      null;
      null;
      null;
      r2910 := (r2643 & r2644 & r2645 & r2646);
      r2911 := rewire_littleendian_2732(r2910);
      null;
      null;
      null;
      null;
      r2913 := (r2647 & r2648 & r2649 & r2650);
      r2914 := rewire_littleendian_2732(r2913);
      null;
      null;
      null;
      null;
      r2916 := (r2651 & r2652 & r2653 & r2654);
      r2917 := rewire_littleendian_2732(r2916);
      null;
      null;
      null;
      null;
      r2919 := (r2655 & r2656 & r2657 & r2658);
      r2920 := rewire_littleendian_2732(r2919);
      null;
      null;
      null;
      null;
      r2922 := (r2659 & r2660 & r2661 & r2662);
      r2923 := rewire_littleendian_2732(r2922);
      null;
      null;
      null;
      null;
      r2925 := (r2663 & r2664 & r2665 & r2666);
      r2926 := rewire_littleendian_2732(r2925);
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      r2928 := (r2881 & r2884 & r2887 & r2890 & r2893 & r2896 & r2899 & r2902 & r2905 & r2908 & r2911 & r2914 & r2917 & r2920 & r2923 & r2926);
      r2601 := r2928;
    end if;
    return r2601;
  end rewire_impwords_2598;
  function rewire_littleendian_2732(r2733 : std_logic_vector) return std_logic_vector
  is
    variable r2878 : std_logic_vector(0 to 31) := (others => '0');
    variable r2877 : std_logic_vector(0 to 15) := (others => '0');
    variable r2876 : std_logic_vector(0 to 15) := (others => '0');
    variable r2830 : std_logic_vector(0 to 15) := (others => '0');
    variable r2829 : std_logic_vector(0 to 7) := (others => '0');
    variable r2828 : std_logic_vector(0 to 7) := (others => '0');
    variable r2749 : std_logic_vector(0 to 31) := (others => '0');
    variable r2748 : std_logic_vector(0 to 15) := (others => '0');
    variable r2747 : std_logic_vector(0 to 15) := (others => '0');
    variable b2745 : boolean := false;
    variable b2744 : boolean := false;
    variable b2743 : boolean := false;
    variable b2742 : boolean := false;
    variable b2741 : boolean := false;
    variable r2740 : std_logic_vector(0 to 7) := (others => '0');
    variable r2739 : std_logic_vector(0 to 7) := (others => '0');
    variable r2738 : std_logic_vector(0 to 7) := (others => '0');
    variable r2737 : std_logic_vector(0 to 7) := (others => '0');
    variable b2736 : boolean := false;
    variable r2735 : std_logic_vector(0 to 31) := (others => '0');
  begin
    b2736 := true;
    r2737 := r2733(0 to 7);
    r2738 := r2733(8 to 15);
    r2739 := r2733(16 to 23);
    r2740 := r2733(24 to 31);
    b2741 := true;
    b2742 := true;
    b2743 := true;
    b2744 := true;
    b2745 := (b2741 AND (b2742 AND (b2743 AND b2744)));
    if b2745 then
      null;
      null;
      r2876 := rewire_w8to16le_2827(r2738,r2737);
      null;
      null;
      r2877 := rewire_w8to16le_2827(r2740,r2739);
      r2878 := rewire_w16tow32le_2746(r2876,r2877);
      r2735 := r2878;
    end if;
    return r2735;
  end rewire_littleendian_2732;
  function rewire_w8to16le_2827(r2828 : std_logic_vector ; r2829 : std_logic_vector) return std_logic_vector
  is
    variable r2875 : std_logic_vector(0 to 15) := (others => '0');
    variable b2873 : boolean := false;
    variable b2872 : boolean := false;
    variable b2871 : boolean := false;
    variable b2870 : boolean := false;
    variable b2869 : boolean := false;
    variable b2868 : boolean := false;
    variable b2867 : boolean := false;
    variable b2866 : boolean := false;
    variable b2865 : boolean := false;
    variable b2864 : boolean := false;
    variable r2863 : std_logic_vector(0 to 0) := (others => '0');
    variable r2862 : std_logic_vector(0 to 0) := (others => '0');
    variable r2861 : std_logic_vector(0 to 0) := (others => '0');
    variable r2860 : std_logic_vector(0 to 0) := (others => '0');
    variable r2859 : std_logic_vector(0 to 0) := (others => '0');
    variable r2858 : std_logic_vector(0 to 0) := (others => '0');
    variable r2857 : std_logic_vector(0 to 0) := (others => '0');
    variable r2856 : std_logic_vector(0 to 0) := (others => '0');
    variable b2855 : boolean := false;
    variable b2854 : boolean := false;
    variable b2853 : boolean := false;
    variable b2852 : boolean := false;
    variable b2851 : boolean := false;
    variable b2850 : boolean := false;
    variable b2849 : boolean := false;
    variable b2848 : boolean := false;
    variable b2847 : boolean := false;
    variable b2846 : boolean := false;
    variable r2845 : std_logic_vector(0 to 0) := (others => '0');
    variable r2844 : std_logic_vector(0 to 0) := (others => '0');
    variable r2843 : std_logic_vector(0 to 0) := (others => '0');
    variable r2842 : std_logic_vector(0 to 0) := (others => '0');
    variable r2841 : std_logic_vector(0 to 0) := (others => '0');
    variable r2840 : std_logic_vector(0 to 0) := (others => '0');
    variable r2839 : std_logic_vector(0 to 0) := (others => '0');
    variable r2838 : std_logic_vector(0 to 0) := (others => '0');
    variable b2837 : boolean := false;
    variable r2836 : std_logic_vector(0 to 7) := (others => '0');
    variable r2835 : std_logic_vector(0 to 7) := (others => '0');
    variable b2834 : boolean := false;
    variable r2833 : std_logic_vector(0 to 15) := (others => '0');
    variable r2832 : std_logic_vector(0 to 15) := (others => '0');
    variable EMPTY : std_logic_vector(0 to -1) := (others => '0');
  begin
    b2834 := true;
    r2835 := r2832(0 to 7);
    r2836 := r2832(8 to 15);
    b2837 := true;
    r2838 := r2835(0 to 0);
    r2839 := r2835(1 to 1);
    r2840 := r2835(2 to 2);
    r2841 := r2835(3 to 3);
    r2842 := r2835(4 to 4);
    r2843 := r2835(5 to 5);
    r2844 := r2835(6 to 6);
    r2845 := r2835(7 to 7);
    b2846 := true;
    b2847 := true;
    b2848 := true;
    b2849 := true;
    b2850 := true;
    b2851 := true;
    b2852 := true;
    b2853 := true;
    b2854 := (b2846 AND (b2847 AND (b2848 AND (b2849 AND (b2850 AND (b2851 AND (b2852 AND b2853)))))));
    b2855 := true;
    r2856 := r2836(0 to 0);
    r2857 := r2836(1 to 1);
    r2858 := r2836(2 to 2);
    r2859 := r2836(3 to 3);
    r2860 := r2836(4 to 4);
    r2861 := r2836(5 to 5);
    r2862 := r2836(6 to 6);
    r2863 := r2836(7 to 7);
    b2864 := true;
    b2865 := true;
    b2866 := true;
    b2867 := true;
    b2868 := true;
    b2869 := true;
    b2870 := true;
    b2871 := true;
    b2872 := (b2864 AND (b2865 AND (b2866 AND (b2867 AND (b2868 AND (b2869 AND (b2870 AND b2871)))))));
    b2873 := (b2854 AND b2872);
    if b2873 then
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      r2875 := (r2856 & r2857 & r2858 & r2859 & r2860 & r2861 & r2862 & r2863 & r2838 & r2839 & r2840 & r2841 & r2842 & r2843 & r2844 & r2845);
      r2833 := r2875;
    end if;
    return r2833;
  end rewire_w8to16le_2827;
  function rewire_w16tow32le_2746(r2747 : std_logic_vector ; r2748 : std_logic_vector) return std_logic_vector
  is
    variable r2826 : std_logic_vector(0 to 31) := (others => '0');
    variable b2824 : boolean := false;
    variable b2823 : boolean := false;
    variable b2822 : boolean := false;
    variable b2821 : boolean := false;
    variable b2820 : boolean := false;
    variable b2819 : boolean := false;
    variable b2818 : boolean := false;
    variable b2817 : boolean := false;
    variable b2816 : boolean := false;
    variable b2815 : boolean := false;
    variable b2814 : boolean := false;
    variable b2813 : boolean := false;
    variable b2812 : boolean := false;
    variable b2811 : boolean := false;
    variable b2810 : boolean := false;
    variable b2809 : boolean := false;
    variable b2808 : boolean := false;
    variable b2807 : boolean := false;
    variable r2806 : std_logic_vector(0 to 0) := (others => '0');
    variable r2805 : std_logic_vector(0 to 0) := (others => '0');
    variable r2804 : std_logic_vector(0 to 0) := (others => '0');
    variable r2803 : std_logic_vector(0 to 0) := (others => '0');
    variable r2802 : std_logic_vector(0 to 0) := (others => '0');
    variable r2801 : std_logic_vector(0 to 0) := (others => '0');
    variable r2800 : std_logic_vector(0 to 0) := (others => '0');
    variable r2799 : std_logic_vector(0 to 0) := (others => '0');
    variable r2798 : std_logic_vector(0 to 0) := (others => '0');
    variable r2797 : std_logic_vector(0 to 0) := (others => '0');
    variable r2796 : std_logic_vector(0 to 0) := (others => '0');
    variable r2795 : std_logic_vector(0 to 0) := (others => '0');
    variable r2794 : std_logic_vector(0 to 0) := (others => '0');
    variable r2793 : std_logic_vector(0 to 0) := (others => '0');
    variable r2792 : std_logic_vector(0 to 0) := (others => '0');
    variable r2791 : std_logic_vector(0 to 0) := (others => '0');
    variable b2790 : boolean := false;
    variable b2789 : boolean := false;
    variable b2788 : boolean := false;
    variable b2787 : boolean := false;
    variable b2786 : boolean := false;
    variable b2785 : boolean := false;
    variable b2784 : boolean := false;
    variable b2783 : boolean := false;
    variable b2782 : boolean := false;
    variable b2781 : boolean := false;
    variable b2780 : boolean := false;
    variable b2779 : boolean := false;
    variable b2778 : boolean := false;
    variable b2777 : boolean := false;
    variable b2776 : boolean := false;
    variable b2775 : boolean := false;
    variable b2774 : boolean := false;
    variable b2773 : boolean := false;
    variable r2772 : std_logic_vector(0 to 0) := (others => '0');
    variable r2771 : std_logic_vector(0 to 0) := (others => '0');
    variable r2770 : std_logic_vector(0 to 0) := (others => '0');
    variable r2769 : std_logic_vector(0 to 0) := (others => '0');
    variable r2768 : std_logic_vector(0 to 0) := (others => '0');
    variable r2767 : std_logic_vector(0 to 0) := (others => '0');
    variable r2766 : std_logic_vector(0 to 0) := (others => '0');
    variable r2765 : std_logic_vector(0 to 0) := (others => '0');
    variable r2764 : std_logic_vector(0 to 0) := (others => '0');
    variable r2763 : std_logic_vector(0 to 0) := (others => '0');
    variable r2762 : std_logic_vector(0 to 0) := (others => '0');
    variable r2761 : std_logic_vector(0 to 0) := (others => '0');
    variable r2760 : std_logic_vector(0 to 0) := (others => '0');
    variable r2759 : std_logic_vector(0 to 0) := (others => '0');
    variable r2758 : std_logic_vector(0 to 0) := (others => '0');
    variable r2757 : std_logic_vector(0 to 0) := (others => '0');
    variable b2756 : boolean := false;
    variable r2755 : std_logic_vector(0 to 15) := (others => '0');
    variable r2754 : std_logic_vector(0 to 15) := (others => '0');
    variable b2753 : boolean := false;
    variable r2752 : std_logic_vector(0 to 31) := (others => '0');
    variable r2751 : std_logic_vector(0 to 31) := (others => '0');
    variable EMPTY : std_logic_vector(0 to -1) := (others => '0');
  begin
    b2753 := true;
    r2754 := r2751(0 to 15);
    r2755 := r2751(16 to 31);
    b2756 := true;
    r2757 := r2754(0 to 0);
    r2758 := r2754(1 to 1);
    r2759 := r2754(2 to 2);
    r2760 := r2754(3 to 3);
    r2761 := r2754(4 to 4);
    r2762 := r2754(5 to 5);
    r2763 := r2754(6 to 6);
    r2764 := r2754(7 to 7);
    r2765 := r2754(8 to 8);
    r2766 := r2754(9 to 9);
    r2767 := r2754(10 to 10);
    r2768 := r2754(11 to 11);
    r2769 := r2754(12 to 12);
    r2770 := r2754(13 to 13);
    r2771 := r2754(14 to 14);
    r2772 := r2754(15 to 15);
    b2773 := true;
    b2774 := true;
    b2775 := true;
    b2776 := true;
    b2777 := true;
    b2778 := true;
    b2779 := true;
    b2780 := true;
    b2781 := true;
    b2782 := true;
    b2783 := true;
    b2784 := true;
    b2785 := true;
    b2786 := true;
    b2787 := true;
    b2788 := true;
    b2789 := (b2773 AND (b2774 AND (b2775 AND (b2776 AND (b2777 AND (b2778 AND (b2779 AND (b2780 AND (b2781 AND (b2782 AND (b2783 AND (b2784 AND (b2785 AND (b2786 AND (b2787 AND b2788)))))))))))))));
    b2790 := true;
    r2791 := r2755(0 to 0);
    r2792 := r2755(1 to 1);
    r2793 := r2755(2 to 2);
    r2794 := r2755(3 to 3);
    r2795 := r2755(4 to 4);
    r2796 := r2755(5 to 5);
    r2797 := r2755(6 to 6);
    r2798 := r2755(7 to 7);
    r2799 := r2755(8 to 8);
    r2800 := r2755(9 to 9);
    r2801 := r2755(10 to 10);
    r2802 := r2755(11 to 11);
    r2803 := r2755(12 to 12);
    r2804 := r2755(13 to 13);
    r2805 := r2755(14 to 14);
    r2806 := r2755(15 to 15);
    b2807 := true;
    b2808 := true;
    b2809 := true;
    b2810 := true;
    b2811 := true;
    b2812 := true;
    b2813 := true;
    b2814 := true;
    b2815 := true;
    b2816 := true;
    b2817 := true;
    b2818 := true;
    b2819 := true;
    b2820 := true;
    b2821 := true;
    b2822 := true;
    b2823 := (b2807 AND (b2808 AND (b2809 AND (b2810 AND (b2811 AND (b2812 AND (b2813 AND (b2814 AND (b2815 AND (b2816 AND (b2817 AND (b2818 AND (b2819 AND (b2820 AND (b2821 AND b2822)))))))))))))));
    b2824 := (b2789 AND b2823);
    if b2824 then
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      r2826 := (r2757 & r2758 & r2759 & r2760 & r2761 & r2762 & r2763 & r2764 & r2765 & r2766 & r2767 & r2768 & r2769 & r2770 & r2771 & r2772 & r2791 & r2792 & r2793 & r2794 & r2795 & r2796 & r2797 & r2798 & r2799 & r2800 & r2801 & r2802 & r2803 & r2804 & r2805 & r2806);
      r2752 := r2826;
    end if;
    return r2752;
  end rewire_w16tow32le_2746;
  function rewire_salsaHashp_1974(r1975 : std_logic_vector) return std_logic_vector
  is
    variable r2597 : std_logic_vector(0 to 511) := (others => '0');
    variable r2596 : std_logic_vector(0 to 31) := (others => '0');
    variable r2595 : std_logic_vector(0 to 31) := (others => '0');
    variable r2594 : std_logic_vector(0 to 31) := (others => '0');
    variable r2593 : std_logic_vector(0 to 31) := (others => '0');
    variable r2592 : std_logic_vector(0 to 31) := (others => '0');
    variable r2591 : std_logic_vector(0 to 31) := (others => '0');
    variable r2590 : std_logic_vector(0 to 31) := (others => '0');
    variable r2589 : std_logic_vector(0 to 31) := (others => '0');
    variable r2588 : std_logic_vector(0 to 31) := (others => '0');
    variable r2587 : std_logic_vector(0 to 31) := (others => '0');
    variable r2586 : std_logic_vector(0 to 31) := (others => '0');
    variable r2585 : std_logic_vector(0 to 31) := (others => '0');
    variable r2584 : std_logic_vector(0 to 31) := (others => '0');
    variable r2583 : std_logic_vector(0 to 31) := (others => '0');
    variable r2582 : std_logic_vector(0 to 31) := (others => '0');
    variable r2581 : std_logic_vector(0 to 31) := (others => '0');
    variable EMPTY : std_logic_vector(0 to -1) := (others => '0');
    variable b2579 : boolean := false;
    variable b2578 : boolean := false;
    variable b2577 : boolean := false;
    variable b2576 : boolean := false;
    variable b2575 : boolean := false;
    variable b2574 : boolean := false;
    variable b2573 : boolean := false;
    variable b2572 : boolean := false;
    variable b2571 : boolean := false;
    variable b2570 : boolean := false;
    variable b2569 : boolean := false;
    variable b2568 : boolean := false;
    variable b2567 : boolean := false;
    variable b2566 : boolean := false;
    variable b2565 : boolean := false;
    variable b2564 : boolean := false;
    variable b2563 : boolean := false;
    variable r2562 : std_logic_vector(0 to 31) := (others => '0');
    variable r2561 : std_logic_vector(0 to 31) := (others => '0');
    variable r2560 : std_logic_vector(0 to 31) := (others => '0');
    variable r2559 : std_logic_vector(0 to 31) := (others => '0');
    variable r2558 : std_logic_vector(0 to 31) := (others => '0');
    variable r2557 : std_logic_vector(0 to 31) := (others => '0');
    variable r2556 : std_logic_vector(0 to 31) := (others => '0');
    variable r2555 : std_logic_vector(0 to 31) := (others => '0');
    variable r2554 : std_logic_vector(0 to 31) := (others => '0');
    variable r2553 : std_logic_vector(0 to 31) := (others => '0');
    variable r2552 : std_logic_vector(0 to 31) := (others => '0');
    variable r2551 : std_logic_vector(0 to 31) := (others => '0');
    variable r2550 : std_logic_vector(0 to 31) := (others => '0');
    variable r2549 : std_logic_vector(0 to 31) := (others => '0');
    variable r2548 : std_logic_vector(0 to 31) := (others => '0');
    variable r2547 : std_logic_vector(0 to 31) := (others => '0');
    variable b2546 : boolean := false;
    variable r2545 : std_logic_vector(0 to 511) := (others => '0');
    variable r2544 : std_logic_vector(0 to 511) := (others => '0');
    variable r2543 : std_logic_vector(0 to 511) := (others => '0');
    variable r2542 : std_logic_vector(0 to 511) := (others => '0');
    variable r2541 : std_logic_vector(0 to 511) := (others => '0');
    variable r2540 : std_logic_vector(0 to 511) := (others => '0');
    variable r2539 : std_logic_vector(0 to 511) := (others => '0');
    variable r2538 : std_logic_vector(0 to 511) := (others => '0');
    variable r2537 : std_logic_vector(0 to 511) := (others => '0');
    variable r2536 : std_logic_vector(0 to 511) := (others => '0');
    variable r2535 : std_logic_vector(0 to 511) := (others => '0');
    variable r2014 : std_logic_vector(0 to 511) := (others => '0');
    variable r2013 : std_logic_vector(0 to 511) := (others => '0');
    variable b2011 : boolean := false;
    variable b2010 : boolean := false;
    variable b2009 : boolean := false;
    variable b2008 : boolean := false;
    variable b2007 : boolean := false;
    variable b2006 : boolean := false;
    variable b2005 : boolean := false;
    variable b2004 : boolean := false;
    variable b2003 : boolean := false;
    variable b2002 : boolean := false;
    variable b2001 : boolean := false;
    variable b2000 : boolean := false;
    variable b1999 : boolean := false;
    variable b1998 : boolean := false;
    variable b1997 : boolean := false;
    variable b1996 : boolean := false;
    variable b1995 : boolean := false;
    variable r1994 : std_logic_vector(0 to 31) := (others => '0');
    variable r1993 : std_logic_vector(0 to 31) := (others => '0');
    variable r1992 : std_logic_vector(0 to 31) := (others => '0');
    variable r1991 : std_logic_vector(0 to 31) := (others => '0');
    variable r1990 : std_logic_vector(0 to 31) := (others => '0');
    variable r1989 : std_logic_vector(0 to 31) := (others => '0');
    variable r1988 : std_logic_vector(0 to 31) := (others => '0');
    variable r1987 : std_logic_vector(0 to 31) := (others => '0');
    variable r1986 : std_logic_vector(0 to 31) := (others => '0');
    variable r1985 : std_logic_vector(0 to 31) := (others => '0');
    variable r1984 : std_logic_vector(0 to 31) := (others => '0');
    variable r1983 : std_logic_vector(0 to 31) := (others => '0');
    variable r1982 : std_logic_vector(0 to 31) := (others => '0');
    variable r1981 : std_logic_vector(0 to 31) := (others => '0');
    variable r1980 : std_logic_vector(0 to 31) := (others => '0');
    variable r1979 : std_logic_vector(0 to 31) := (others => '0');
    variable b1978 : boolean := false;
    variable r1977 : std_logic_vector(0 to 511) := (others => '0');
  begin
    b1978 := true;
    r1979 := r1975(0 to 31);
    r1980 := r1975(32 to 63);
    r1981 := r1975(64 to 95);
    r1982 := r1975(96 to 127);
    r1983 := r1975(128 to 159);
    r1984 := r1975(160 to 191);
    r1985 := r1975(192 to 223);
    r1986 := r1975(224 to 255);
    r1987 := r1975(256 to 287);
    r1988 := r1975(288 to 319);
    r1989 := r1975(320 to 351);
    r1990 := r1975(352 to 383);
    r1991 := r1975(384 to 415);
    r1992 := r1975(416 to 447);
    r1993 := r1975(448 to 479);
    r1994 := r1975(480 to 511);
    b1995 := true;
    b1996 := true;
    b1997 := true;
    b1998 := true;
    b1999 := true;
    b2000 := true;
    b2001 := true;
    b2002 := true;
    b2003 := true;
    b2004 := true;
    b2005 := true;
    b2006 := true;
    b2007 := true;
    b2008 := true;
    b2009 := true;
    b2010 := true;
    b2011 := (b1995 AND (b1996 AND (b1997 AND (b1998 AND (b1999 AND (b2000 AND (b2001 AND (b2002 AND (b2003 AND (b2004 AND (b2005 AND (b2006 AND (b2007 AND (b2008 AND (b2009 AND b2010)))))))))))))));
    if b2011 then
      b2546 := true;
      r2547 := r2544(0 to 31);
      r2548 := r2544(32 to 63);
      r2549 := r2544(64 to 95);
      r2550 := r2544(96 to 127);
      r2551 := r2544(128 to 159);
      r2552 := r2544(160 to 191);
      r2553 := r2544(192 to 223);
      r2554 := r2544(224 to 255);
      r2555 := r2544(256 to 287);
      r2556 := r2544(288 to 319);
      r2557 := r2544(320 to 351);
      r2558 := r2544(352 to 383);
      r2559 := r2544(384 to 415);
      r2560 := r2544(416 to 447);
      r2561 := r2544(448 to 479);
      r2562 := r2544(480 to 511);
      b2563 := true;
      b2564 := true;
      b2565 := true;
      b2566 := true;
      b2567 := true;
      b2568 := true;
      b2569 := true;
      b2570 := true;
      b2571 := true;
      b2572 := true;
      b2573 := true;
      b2574 := true;
      b2575 := true;
      b2576 := true;
      b2577 := true;
      b2578 := true;
      b2579 := (b2563 AND (b2564 AND (b2565 AND (b2566 AND (b2567 AND (b2568 AND (b2569 AND (b2570 AND (b2571 AND (b2572 AND (b2573 AND (b2574 AND (b2575 AND (b2576 AND (b2577 AND b2578)))))))))))))));
      if b2579 then
        null;
        null;
        r2581 := add32(r2547,r1979);
        null;
        null;
        r2582 := add32(r2548,r1980);
        null;
        null;
        r2583 := add32(r2549,r1981);
        null;
        null;
        r2584 := add32(r2550,r1982);
        null;
        null;
        r2585 := add32(r2551,r1983);
        null;
        null;
        r2586 := add32(r2552,r1984);
        null;
        null;
        r2587 := add32(r2553,r1985);
        null;
        null;
        r2588 := add32(r2554,r1986);
        null;
        null;
        r2589 := add32(r2555,r1987);
        null;
        null;
        r2590 := add32(r2556,r1988);
        null;
        null;
        r2591 := add32(r2557,r1989);
        null;
        null;
        r2592 := add32(r2558,r1990);
        null;
        null;
        r2593 := add32(r2559,r1991);
        null;
        null;
        r2594 := add32(r2560,r1992);
        null;
        null;
        r2595 := add32(r2561,r1993);
        null;
        null;
        r2596 := add32(r2562,r1994);
        r2597 := (r2581 & r2582 & r2583 & r2584 & r2585 & r2586 & r2587 & r2588 & r2589 & r2590 & r2591 & r2592 & r2593 & r2594 & r2595 & r2596);
        r2545 := r2597;
      end if;
      r1977 := r2545;
    end if;
    return r1977;
  end rewire_salsaHashp_1974;
  function rewire_doubleRound_2012(r2013 : std_logic_vector) return std_logic_vector
  is
    variable r2534 : std_logic_vector(0 to 511) := (others => '0');
    variable r2533 : std_logic_vector(0 to 511) := (others => '0');
    variable r2434 : std_logic_vector(0 to 511) := (others => '0');
    variable r2433 : std_logic_vector(0 to 511) := (others => '0');
    variable r2017 : std_logic_vector(0 to 511) := (others => '0');
    variable r2016 : std_logic_vector(0 to 511) := (others => '0');
  begin
    null;
    r2533 := rewire_columnRound_2432(r2013);
    r2534 := rewire_rowRound_2015(r2533);
    return r2534;
  end rewire_doubleRound_2012;
  function rewire_columnRound_2432(r2433 : std_logic_vector) return std_logic_vector
  is
    variable r2532 : std_logic_vector(0 to 511) := (others => '0');
    variable b2530 : boolean := false;
    variable b2529 : boolean := false;
    variable b2528 : boolean := false;
    variable b2527 : boolean := false;
    variable b2526 : boolean := false;
    variable b2525 : boolean := false;
    variable r2524 : std_logic_vector(0 to 31) := (others => '0');
    variable r2523 : std_logic_vector(0 to 31) := (others => '0');
    variable r2522 : std_logic_vector(0 to 31) := (others => '0');
    variable r2521 : std_logic_vector(0 to 31) := (others => '0');
    variable b2520 : boolean := false;
    variable b2519 : boolean := false;
    variable b2518 : boolean := false;
    variable b2517 : boolean := false;
    variable b2516 : boolean := false;
    variable b2515 : boolean := false;
    variable r2514 : std_logic_vector(0 to 31) := (others => '0');
    variable r2513 : std_logic_vector(0 to 31) := (others => '0');
    variable r2512 : std_logic_vector(0 to 31) := (others => '0');
    variable r2511 : std_logic_vector(0 to 31) := (others => '0');
    variable b2510 : boolean := false;
    variable b2509 : boolean := false;
    variable b2508 : boolean := false;
    variable b2507 : boolean := false;
    variable b2506 : boolean := false;
    variable b2505 : boolean := false;
    variable r2504 : std_logic_vector(0 to 31) := (others => '0');
    variable r2503 : std_logic_vector(0 to 31) := (others => '0');
    variable r2502 : std_logic_vector(0 to 31) := (others => '0');
    variable r2501 : std_logic_vector(0 to 31) := (others => '0');
    variable b2500 : boolean := false;
    variable b2499 : boolean := false;
    variable b2498 : boolean := false;
    variable b2497 : boolean := false;
    variable b2496 : boolean := false;
    variable b2495 : boolean := false;
    variable r2494 : std_logic_vector(0 to 31) := (others => '0');
    variable r2493 : std_logic_vector(0 to 31) := (others => '0');
    variable r2492 : std_logic_vector(0 to 31) := (others => '0');
    variable r2491 : std_logic_vector(0 to 31) := (others => '0');
    variable b2490 : boolean := false;
    variable r2489 : std_logic_vector(0 to 127) := (others => '0');
    variable r2488 : std_logic_vector(0 to 127) := (others => '0');
    variable r2487 : std_logic_vector(0 to 127) := (others => '0');
    variable r2486 : std_logic_vector(0 to 127) := (others => '0');
    variable b2485 : boolean := false;
    variable r2484 : std_logic_vector(0 to 511) := (others => '0');
    variable r2483 : std_logic_vector(0 to 511) := (others => '0');
    variable r2481 : std_logic_vector(0 to 127) := (others => '0');
    variable r2480 : std_logic_vector(0 to 127) := (others => '0');
    variable r2478 : std_logic_vector(0 to 127) := (others => '0');
    variable r2477 : std_logic_vector(0 to 127) := (others => '0');
    variable r2475 : std_logic_vector(0 to 127) := (others => '0');
    variable r2474 : std_logic_vector(0 to 127) := (others => '0');
    variable r2472 : std_logic_vector(0 to 127) := (others => '0');
    variable r2471 : std_logic_vector(0 to 127) := (others => '0');
    variable EMPTY : std_logic_vector(0 to -1) := (others => '0');
    variable b2469 : boolean := false;
    variable b2468 : boolean := false;
    variable b2467 : boolean := false;
    variable b2466 : boolean := false;
    variable b2465 : boolean := false;
    variable b2464 : boolean := false;
    variable b2463 : boolean := false;
    variable b2462 : boolean := false;
    variable b2461 : boolean := false;
    variable b2460 : boolean := false;
    variable b2459 : boolean := false;
    variable b2458 : boolean := false;
    variable b2457 : boolean := false;
    variable b2456 : boolean := false;
    variable b2455 : boolean := false;
    variable b2454 : boolean := false;
    variable b2453 : boolean := false;
    variable r2452 : std_logic_vector(0 to 31) := (others => '0');
    variable r2451 : std_logic_vector(0 to 31) := (others => '0');
    variable r2450 : std_logic_vector(0 to 31) := (others => '0');
    variable r2449 : std_logic_vector(0 to 31) := (others => '0');
    variable r2448 : std_logic_vector(0 to 31) := (others => '0');
    variable r2447 : std_logic_vector(0 to 31) := (others => '0');
    variable r2446 : std_logic_vector(0 to 31) := (others => '0');
    variable r2445 : std_logic_vector(0 to 31) := (others => '0');
    variable r2444 : std_logic_vector(0 to 31) := (others => '0');
    variable r2443 : std_logic_vector(0 to 31) := (others => '0');
    variable r2442 : std_logic_vector(0 to 31) := (others => '0');
    variable r2441 : std_logic_vector(0 to 31) := (others => '0');
    variable r2440 : std_logic_vector(0 to 31) := (others => '0');
    variable r2439 : std_logic_vector(0 to 31) := (others => '0');
    variable r2438 : std_logic_vector(0 to 31) := (others => '0');
    variable r2437 : std_logic_vector(0 to 31) := (others => '0');
    variable b2436 : boolean := false;
    variable r2435 : std_logic_vector(0 to 511) := (others => '0');
  begin
    b2436 := true;
    r2437 := r2433(0 to 31);
    r2438 := r2433(32 to 63);
    r2439 := r2433(64 to 95);
    r2440 := r2433(96 to 127);
    r2441 := r2433(128 to 159);
    r2442 := r2433(160 to 191);
    r2443 := r2433(192 to 223);
    r2444 := r2433(224 to 255);
    r2445 := r2433(256 to 287);
    r2446 := r2433(288 to 319);
    r2447 := r2433(320 to 351);
    r2448 := r2433(352 to 383);
    r2449 := r2433(384 to 415);
    r2450 := r2433(416 to 447);
    r2451 := r2433(448 to 479);
    r2452 := r2433(480 to 511);
    b2453 := true;
    b2454 := true;
    b2455 := true;
    b2456 := true;
    b2457 := true;
    b2458 := true;
    b2459 := true;
    b2460 := true;
    b2461 := true;
    b2462 := true;
    b2463 := true;
    b2464 := true;
    b2465 := true;
    b2466 := true;
    b2467 := true;
    b2468 := true;
    b2469 := (b2453 AND (b2454 AND (b2455 AND (b2456 AND (b2457 AND (b2458 AND (b2459 AND (b2460 AND (b2461 AND (b2462 AND (b2463 AND (b2464 AND (b2465 AND (b2466 AND (b2467 AND b2468)))))))))))))));
    if b2469 then
      null;
      null;
      null;
      null;
      r2471 := (r2437 & r2441 & r2445 & r2449);
      r2472 := rewire_quarterRound_2053(r2471);
      null;
      null;
      null;
      null;
      r2474 := (r2442 & r2446 & r2450 & r2438);
      r2475 := rewire_quarterRound_2053(r2474);
      null;
      null;
      null;
      null;
      r2477 := (r2447 & r2451 & r2439 & r2443);
      r2478 := rewire_quarterRound_2053(r2477);
      null;
      null;
      null;
      null;
      r2480 := (r2452 & r2440 & r2444 & r2448);
      r2481 := rewire_quarterRound_2053(r2480);
      b2485 := true;
      r2486 := r2483(0 to 127);
      r2487 := r2483(128 to 255);
      r2488 := r2483(256 to 383);
      r2489 := r2483(384 to 511);
      b2490 := true;
      r2491 := r2486(0 to 31);
      r2492 := r2486(32 to 63);
      r2493 := r2486(64 to 95);
      r2494 := r2486(96 to 127);
      b2495 := true;
      b2496 := true;
      b2497 := true;
      b2498 := true;
      b2499 := (b2495 AND (b2496 AND (b2497 AND b2498)));
      b2500 := true;
      r2501 := r2487(0 to 31);
      r2502 := r2487(32 to 63);
      r2503 := r2487(64 to 95);
      r2504 := r2487(96 to 127);
      b2505 := true;
      b2506 := true;
      b2507 := true;
      b2508 := true;
      b2509 := (b2505 AND (b2506 AND (b2507 AND b2508)));
      b2510 := true;
      r2511 := r2488(0 to 31);
      r2512 := r2488(32 to 63);
      r2513 := r2488(64 to 95);
      r2514 := r2488(96 to 127);
      b2515 := true;
      b2516 := true;
      b2517 := true;
      b2518 := true;
      b2519 := (b2515 AND (b2516 AND (b2517 AND b2518)));
      b2520 := true;
      r2521 := r2489(0 to 31);
      r2522 := r2489(32 to 63);
      r2523 := r2489(64 to 95);
      r2524 := r2489(96 to 127);
      b2525 := true;
      b2526 := true;
      b2527 := true;
      b2528 := true;
      b2529 := (b2525 AND (b2526 AND (b2527 AND b2528)));
      b2530 := (b2499 AND (b2509 AND (b2519 AND b2529)));
      if b2530 then
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        r2532 := (r2491 & r2504 & r2513 & r2522 & r2492 & r2501 & r2514 & r2523 & r2493 & r2502 & r2511 & r2524 & r2494 & r2503 & r2512 & r2521);
        r2484 := r2532;
      end if;
      r2435 := r2484;
    end if;
    return r2435;
  end rewire_columnRound_2432;
  function rewire_rowRound_2015(r2016 : std_logic_vector) return std_logic_vector
  is
    variable r2431 : std_logic_vector(0 to 511) := (others => '0');
    variable b2429 : boolean := false;
    variable b2428 : boolean := false;
    variable b2427 : boolean := false;
    variable b2426 : boolean := false;
    variable b2425 : boolean := false;
    variable b2424 : boolean := false;
    variable r2423 : std_logic_vector(0 to 31) := (others => '0');
    variable r2422 : std_logic_vector(0 to 31) := (others => '0');
    variable r2421 : std_logic_vector(0 to 31) := (others => '0');
    variable r2420 : std_logic_vector(0 to 31) := (others => '0');
    variable b2419 : boolean := false;
    variable b2418 : boolean := false;
    variable b2417 : boolean := false;
    variable b2416 : boolean := false;
    variable b2415 : boolean := false;
    variable b2414 : boolean := false;
    variable r2413 : std_logic_vector(0 to 31) := (others => '0');
    variable r2412 : std_logic_vector(0 to 31) := (others => '0');
    variable r2411 : std_logic_vector(0 to 31) := (others => '0');
    variable r2410 : std_logic_vector(0 to 31) := (others => '0');
    variable b2409 : boolean := false;
    variable b2408 : boolean := false;
    variable b2407 : boolean := false;
    variable b2406 : boolean := false;
    variable b2405 : boolean := false;
    variable b2404 : boolean := false;
    variable r2403 : std_logic_vector(0 to 31) := (others => '0');
    variable r2402 : std_logic_vector(0 to 31) := (others => '0');
    variable r2401 : std_logic_vector(0 to 31) := (others => '0');
    variable r2400 : std_logic_vector(0 to 31) := (others => '0');
    variable b2399 : boolean := false;
    variable b2398 : boolean := false;
    variable b2397 : boolean := false;
    variable b2396 : boolean := false;
    variable b2395 : boolean := false;
    variable b2394 : boolean := false;
    variable r2393 : std_logic_vector(0 to 31) := (others => '0');
    variable r2392 : std_logic_vector(0 to 31) := (others => '0');
    variable r2391 : std_logic_vector(0 to 31) := (others => '0');
    variable r2390 : std_logic_vector(0 to 31) := (others => '0');
    variable b2389 : boolean := false;
    variable r2388 : std_logic_vector(0 to 127) := (others => '0');
    variable r2387 : std_logic_vector(0 to 127) := (others => '0');
    variable r2386 : std_logic_vector(0 to 127) := (others => '0');
    variable r2385 : std_logic_vector(0 to 127) := (others => '0');
    variable b2384 : boolean := false;
    variable r2383 : std_logic_vector(0 to 511) := (others => '0');
    variable r2382 : std_logic_vector(0 to 511) := (others => '0');
    variable r2380 : std_logic_vector(0 to 127) := (others => '0');
    variable r2379 : std_logic_vector(0 to 127) := (others => '0');
    variable r2377 : std_logic_vector(0 to 127) := (others => '0');
    variable r2376 : std_logic_vector(0 to 127) := (others => '0');
    variable r2374 : std_logic_vector(0 to 127) := (others => '0');
    variable r2373 : std_logic_vector(0 to 127) := (others => '0');
    variable r2371 : std_logic_vector(0 to 127) := (others => '0');
    variable r2370 : std_logic_vector(0 to 127) := (others => '0');
    variable EMPTY : std_logic_vector(0 to -1) := (others => '0');
    variable r2055 : std_logic_vector(0 to 127) := (others => '0');
    variable r2054 : std_logic_vector(0 to 127) := (others => '0');
    variable b2052 : boolean := false;
    variable b2051 : boolean := false;
    variable b2050 : boolean := false;
    variable b2049 : boolean := false;
    variable b2048 : boolean := false;
    variable b2047 : boolean := false;
    variable b2046 : boolean := false;
    variable b2045 : boolean := false;
    variable b2044 : boolean := false;
    variable b2043 : boolean := false;
    variable b2042 : boolean := false;
    variable b2041 : boolean := false;
    variable b2040 : boolean := false;
    variable b2039 : boolean := false;
    variable b2038 : boolean := false;
    variable b2037 : boolean := false;
    variable b2036 : boolean := false;
    variable r2035 : std_logic_vector(0 to 31) := (others => '0');
    variable r2034 : std_logic_vector(0 to 31) := (others => '0');
    variable r2033 : std_logic_vector(0 to 31) := (others => '0');
    variable r2032 : std_logic_vector(0 to 31) := (others => '0');
    variable r2031 : std_logic_vector(0 to 31) := (others => '0');
    variable r2030 : std_logic_vector(0 to 31) := (others => '0');
    variable r2029 : std_logic_vector(0 to 31) := (others => '0');
    variable r2028 : std_logic_vector(0 to 31) := (others => '0');
    variable r2027 : std_logic_vector(0 to 31) := (others => '0');
    variable r2026 : std_logic_vector(0 to 31) := (others => '0');
    variable r2025 : std_logic_vector(0 to 31) := (others => '0');
    variable r2024 : std_logic_vector(0 to 31) := (others => '0');
    variable r2023 : std_logic_vector(0 to 31) := (others => '0');
    variable r2022 : std_logic_vector(0 to 31) := (others => '0');
    variable r2021 : std_logic_vector(0 to 31) := (others => '0');
    variable r2020 : std_logic_vector(0 to 31) := (others => '0');
    variable b2019 : boolean := false;
    variable r2018 : std_logic_vector(0 to 511) := (others => '0');
  begin
    b2019 := true;
    r2020 := r2016(0 to 31);
    r2021 := r2016(32 to 63);
    r2022 := r2016(64 to 95);
    r2023 := r2016(96 to 127);
    r2024 := r2016(128 to 159);
    r2025 := r2016(160 to 191);
    r2026 := r2016(192 to 223);
    r2027 := r2016(224 to 255);
    r2028 := r2016(256 to 287);
    r2029 := r2016(288 to 319);
    r2030 := r2016(320 to 351);
    r2031 := r2016(352 to 383);
    r2032 := r2016(384 to 415);
    r2033 := r2016(416 to 447);
    r2034 := r2016(448 to 479);
    r2035 := r2016(480 to 511);
    b2036 := true;
    b2037 := true;
    b2038 := true;
    b2039 := true;
    b2040 := true;
    b2041 := true;
    b2042 := true;
    b2043 := true;
    b2044 := true;
    b2045 := true;
    b2046 := true;
    b2047 := true;
    b2048 := true;
    b2049 := true;
    b2050 := true;
    b2051 := true;
    b2052 := (b2036 AND (b2037 AND (b2038 AND (b2039 AND (b2040 AND (b2041 AND (b2042 AND (b2043 AND (b2044 AND (b2045 AND (b2046 AND (b2047 AND (b2048 AND (b2049 AND (b2050 AND b2051)))))))))))))));
    if b2052 then
      null;
      null;
      null;
      null;
      r2370 := (r2020 & r2021 & r2022 & r2023);
      r2371 := rewire_quarterRound_2053(r2370);
      null;
      null;
      null;
      null;
      r2373 := (r2025 & r2026 & r2027 & r2024);
      r2374 := rewire_quarterRound_2053(r2373);
      null;
      null;
      null;
      null;
      r2376 := (r2030 & r2031 & r2028 & r2029);
      r2377 := rewire_quarterRound_2053(r2376);
      null;
      null;
      null;
      null;
      r2379 := (r2035 & r2032 & r2033 & r2034);
      r2380 := rewire_quarterRound_2053(r2379);
      b2384 := true;
      r2385 := r2382(0 to 127);
      r2386 := r2382(128 to 255);
      r2387 := r2382(256 to 383);
      r2388 := r2382(384 to 511);
      b2389 := true;
      r2390 := r2385(0 to 31);
      r2391 := r2385(32 to 63);
      r2392 := r2385(64 to 95);
      r2393 := r2385(96 to 127);
      b2394 := true;
      b2395 := true;
      b2396 := true;
      b2397 := true;
      b2398 := (b2394 AND (b2395 AND (b2396 AND b2397)));
      b2399 := true;
      r2400 := r2386(0 to 31);
      r2401 := r2386(32 to 63);
      r2402 := r2386(64 to 95);
      r2403 := r2386(96 to 127);
      b2404 := true;
      b2405 := true;
      b2406 := true;
      b2407 := true;
      b2408 := (b2404 AND (b2405 AND (b2406 AND b2407)));
      b2409 := true;
      r2410 := r2387(0 to 31);
      r2411 := r2387(32 to 63);
      r2412 := r2387(64 to 95);
      r2413 := r2387(96 to 127);
      b2414 := true;
      b2415 := true;
      b2416 := true;
      b2417 := true;
      b2418 := (b2414 AND (b2415 AND (b2416 AND b2417)));
      b2419 := true;
      r2420 := r2388(0 to 31);
      r2421 := r2388(32 to 63);
      r2422 := r2388(64 to 95);
      r2423 := r2388(96 to 127);
      b2424 := true;
      b2425 := true;
      b2426 := true;
      b2427 := true;
      b2428 := (b2424 AND (b2425 AND (b2426 AND b2427)));
      b2429 := (b2398 AND (b2408 AND (b2418 AND b2428)));
      if b2429 then
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        r2431 := (r2390 & r2391 & r2392 & r2393 & r2403 & r2400 & r2401 & r2402 & r2412 & r2413 & r2410 & r2411 & r2421 & r2422 & r2423 & r2420);
        r2383 := r2431;
      end if;
      r2018 := r2383;
    end if;
    return r2018;
  end rewire_rowRound_2015;
  function rewire_quarterRound_2053(r2054 : std_logic_vector) return std_logic_vector
  is
    variable r2368 : std_logic_vector(0 to 127) := (others => '0');
    variable EMPTY : std_logic_vector(0 to -1) := (others => '0');
    variable r2366 : std_logic_vector(0 to 31) := (others => '0');
    variable r2365 : std_logic_vector(0 to 31) := (others => '0');
    variable r2364 : std_logic_vector(0 to 31) := (others => '0');
    variable r2294 : std_logic_vector(0 to 31) := (others => '0');
    variable r2293 : std_logic_vector(0 to 31) := (others => '0');
    variable r2291 : std_logic_vector(0 to 31) := (others => '0');
    variable r2290 : std_logic_vector(0 to 31) := (others => '0');
    variable r2289 : std_logic_vector(0 to 31) := (others => '0');
    variable r2219 : std_logic_vector(0 to 31) := (others => '0');
    variable r2218 : std_logic_vector(0 to 31) := (others => '0');
    variable r2216 : std_logic_vector(0 to 31) := (others => '0');
    variable r2215 : std_logic_vector(0 to 31) := (others => '0');
    variable r2214 : std_logic_vector(0 to 31) := (others => '0');
    variable r2144 : std_logic_vector(0 to 31) := (others => '0');
    variable r2143 : std_logic_vector(0 to 31) := (others => '0');
    variable r2141 : std_logic_vector(0 to 31) := (others => '0');
    variable r2140 : std_logic_vector(0 to 31) := (others => '0');
    variable r2139 : std_logic_vector(0 to 31) := (others => '0');
    variable r2069 : std_logic_vector(0 to 31) := (others => '0');
    variable r2068 : std_logic_vector(0 to 31) := (others => '0');
    variable b2066 : boolean := false;
    variable b2065 : boolean := false;
    variable b2064 : boolean := false;
    variable b2063 : boolean := false;
    variable b2062 : boolean := false;
    variable r2061 : std_logic_vector(0 to 31) := (others => '0');
    variable r2060 : std_logic_vector(0 to 31) := (others => '0');
    variable r2059 : std_logic_vector(0 to 31) := (others => '0');
    variable r2058 : std_logic_vector(0 to 31) := (others => '0');
    variable b2057 : boolean := false;
    variable r2056 : std_logic_vector(0 to 127) := (others => '0');
  begin
    b2057 := true;
    r2058 := r2054(0 to 31);
    r2059 := r2054(32 to 63);
    r2060 := r2054(64 to 95);
    r2061 := r2054(96 to 127);
    b2062 := true;
    b2063 := true;
    b2064 := true;
    b2065 := true;
    b2066 := (b2062 AND (b2063 AND (b2064 AND b2065)));
    if b2066 then
      null;
      null;
      null;
      r2139 := add32(r2058,r2061);
      r2140 := rewire_rot7_2067(r2139);
      r2141 := xor32(r2059,r2140);
      null;
      null;
      null;
      r2214 := add32(r2141,r2058);
      r2215 := rewire_rot9_2142(r2214);
      r2216 := xor32(r2060,r2215);
      null;
      null;
      null;
      r2289 := add32(r2216,r2141);
      r2290 := rewire_rot13_2217(r2289);
      r2291 := xor32(r2061,r2290);
      null;
      null;
      null;
      r2364 := add32(r2291,r2216);
      r2365 := rewire_rot18_2292(r2364);
      r2366 := xor32(r2058,r2365);
      null;
      null;
      null;
      null;
      r2368 := (r2366 & r2141 & r2216 & r2291);
      r2056 := r2368;
    end if;
    return r2056;
  end rewire_quarterRound_2053;
  function rewire_rot18_2292(r2293 : std_logic_vector) return std_logic_vector
  is
    variable r2363 : std_logic_vector(0 to 31) := (others => '0');
    variable EMPTY : std_logic_vector(0 to -1) := (others => '0');
    variable b2361 : boolean := false;
    variable b2360 : boolean := false;
    variable b2359 : boolean := false;
    variable b2358 : boolean := false;
    variable b2357 : boolean := false;
    variable b2356 : boolean := false;
    variable b2355 : boolean := false;
    variable b2354 : boolean := false;
    variable b2353 : boolean := false;
    variable b2352 : boolean := false;
    variable b2351 : boolean := false;
    variable b2350 : boolean := false;
    variable b2349 : boolean := false;
    variable b2348 : boolean := false;
    variable b2347 : boolean := false;
    variable b2346 : boolean := false;
    variable b2345 : boolean := false;
    variable b2344 : boolean := false;
    variable b2343 : boolean := false;
    variable b2342 : boolean := false;
    variable b2341 : boolean := false;
    variable b2340 : boolean := false;
    variable b2339 : boolean := false;
    variable b2338 : boolean := false;
    variable b2337 : boolean := false;
    variable b2336 : boolean := false;
    variable b2335 : boolean := false;
    variable b2334 : boolean := false;
    variable b2333 : boolean := false;
    variable b2332 : boolean := false;
    variable b2331 : boolean := false;
    variable b2330 : boolean := false;
    variable b2329 : boolean := false;
    variable r2328 : std_logic_vector(0 to 0) := (others => '0');
    variable r2327 : std_logic_vector(0 to 0) := (others => '0');
    variable r2326 : std_logic_vector(0 to 0) := (others => '0');
    variable r2325 : std_logic_vector(0 to 0) := (others => '0');
    variable r2324 : std_logic_vector(0 to 0) := (others => '0');
    variable r2323 : std_logic_vector(0 to 0) := (others => '0');
    variable r2322 : std_logic_vector(0 to 0) := (others => '0');
    variable r2321 : std_logic_vector(0 to 0) := (others => '0');
    variable r2320 : std_logic_vector(0 to 0) := (others => '0');
    variable r2319 : std_logic_vector(0 to 0) := (others => '0');
    variable r2318 : std_logic_vector(0 to 0) := (others => '0');
    variable r2317 : std_logic_vector(0 to 0) := (others => '0');
    variable r2316 : std_logic_vector(0 to 0) := (others => '0');
    variable r2315 : std_logic_vector(0 to 0) := (others => '0');
    variable r2314 : std_logic_vector(0 to 0) := (others => '0');
    variable r2313 : std_logic_vector(0 to 0) := (others => '0');
    variable r2312 : std_logic_vector(0 to 0) := (others => '0');
    variable r2311 : std_logic_vector(0 to 0) := (others => '0');
    variable r2310 : std_logic_vector(0 to 0) := (others => '0');
    variable r2309 : std_logic_vector(0 to 0) := (others => '0');
    variable r2308 : std_logic_vector(0 to 0) := (others => '0');
    variable r2307 : std_logic_vector(0 to 0) := (others => '0');
    variable r2306 : std_logic_vector(0 to 0) := (others => '0');
    variable r2305 : std_logic_vector(0 to 0) := (others => '0');
    variable r2304 : std_logic_vector(0 to 0) := (others => '0');
    variable r2303 : std_logic_vector(0 to 0) := (others => '0');
    variable r2302 : std_logic_vector(0 to 0) := (others => '0');
    variable r2301 : std_logic_vector(0 to 0) := (others => '0');
    variable r2300 : std_logic_vector(0 to 0) := (others => '0');
    variable r2299 : std_logic_vector(0 to 0) := (others => '0');
    variable r2298 : std_logic_vector(0 to 0) := (others => '0');
    variable r2297 : std_logic_vector(0 to 0) := (others => '0');
    variable b2296 : boolean := false;
    variable r2295 : std_logic_vector(0 to 31) := (others => '0');
  begin
    b2296 := true;
    r2297 := r2293(0 to 0);
    r2298 := r2293(1 to 1);
    r2299 := r2293(2 to 2);
    r2300 := r2293(3 to 3);
    r2301 := r2293(4 to 4);
    r2302 := r2293(5 to 5);
    r2303 := r2293(6 to 6);
    r2304 := r2293(7 to 7);
    r2305 := r2293(8 to 8);
    r2306 := r2293(9 to 9);
    r2307 := r2293(10 to 10);
    r2308 := r2293(11 to 11);
    r2309 := r2293(12 to 12);
    r2310 := r2293(13 to 13);
    r2311 := r2293(14 to 14);
    r2312 := r2293(15 to 15);
    r2313 := r2293(16 to 16);
    r2314 := r2293(17 to 17);
    r2315 := r2293(18 to 18);
    r2316 := r2293(19 to 19);
    r2317 := r2293(20 to 20);
    r2318 := r2293(21 to 21);
    r2319 := r2293(22 to 22);
    r2320 := r2293(23 to 23);
    r2321 := r2293(24 to 24);
    r2322 := r2293(25 to 25);
    r2323 := r2293(26 to 26);
    r2324 := r2293(27 to 27);
    r2325 := r2293(28 to 28);
    r2326 := r2293(29 to 29);
    r2327 := r2293(30 to 30);
    r2328 := r2293(31 to 31);
    b2329 := true;
    b2330 := true;
    b2331 := true;
    b2332 := true;
    b2333 := true;
    b2334 := true;
    b2335 := true;
    b2336 := true;
    b2337 := true;
    b2338 := true;
    b2339 := true;
    b2340 := true;
    b2341 := true;
    b2342 := true;
    b2343 := true;
    b2344 := true;
    b2345 := true;
    b2346 := true;
    b2347 := true;
    b2348 := true;
    b2349 := true;
    b2350 := true;
    b2351 := true;
    b2352 := true;
    b2353 := true;
    b2354 := true;
    b2355 := true;
    b2356 := true;
    b2357 := true;
    b2358 := true;
    b2359 := true;
    b2360 := true;
    b2361 := (b2329 AND (b2330 AND (b2331 AND (b2332 AND (b2333 AND (b2334 AND (b2335 AND (b2336 AND (b2337 AND (b2338 AND (b2339 AND (b2340 AND (b2341 AND (b2342 AND (b2343 AND (b2344 AND (b2345 AND (b2346 AND (b2347 AND (b2348 AND (b2349 AND (b2350 AND (b2351 AND (b2352 AND (b2353 AND (b2354 AND (b2355 AND (b2356 AND (b2357 AND (b2358 AND (b2359 AND b2360)))))))))))))))))))))))))))))));
    if b2361 then
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      r2363 := (r2311 & r2312 & r2313 & r2314 & r2315 & r2316 & r2317 & r2318 & r2319 & r2320 & r2321 & r2322 & r2323 & r2324 & r2325 & r2326 & r2327 & r2328 & r2297 & r2298 & r2299 & r2300 & r2301 & r2302 & r2303 & r2304 & r2305 & r2306 & r2307 & r2308 & r2309 & r2310);
      r2295 := r2363;
    end if;
    return r2295;
  end rewire_rot18_2292;
  function rewire_rot13_2217(r2218 : std_logic_vector) return std_logic_vector
  is
    variable r2288 : std_logic_vector(0 to 31) := (others => '0');
    variable EMPTY : std_logic_vector(0 to -1) := (others => '0');
    variable b2286 : boolean := false;
    variable b2285 : boolean := false;
    variable b2284 : boolean := false;
    variable b2283 : boolean := false;
    variable b2282 : boolean := false;
    variable b2281 : boolean := false;
    variable b2280 : boolean := false;
    variable b2279 : boolean := false;
    variable b2278 : boolean := false;
    variable b2277 : boolean := false;
    variable b2276 : boolean := false;
    variable b2275 : boolean := false;
    variable b2274 : boolean := false;
    variable b2273 : boolean := false;
    variable b2272 : boolean := false;
    variable b2271 : boolean := false;
    variable b2270 : boolean := false;
    variable b2269 : boolean := false;
    variable b2268 : boolean := false;
    variable b2267 : boolean := false;
    variable b2266 : boolean := false;
    variable b2265 : boolean := false;
    variable b2264 : boolean := false;
    variable b2263 : boolean := false;
    variable b2262 : boolean := false;
    variable b2261 : boolean := false;
    variable b2260 : boolean := false;
    variable b2259 : boolean := false;
    variable b2258 : boolean := false;
    variable b2257 : boolean := false;
    variable b2256 : boolean := false;
    variable b2255 : boolean := false;
    variable b2254 : boolean := false;
    variable r2253 : std_logic_vector(0 to 0) := (others => '0');
    variable r2252 : std_logic_vector(0 to 0) := (others => '0');
    variable r2251 : std_logic_vector(0 to 0) := (others => '0');
    variable r2250 : std_logic_vector(0 to 0) := (others => '0');
    variable r2249 : std_logic_vector(0 to 0) := (others => '0');
    variable r2248 : std_logic_vector(0 to 0) := (others => '0');
    variable r2247 : std_logic_vector(0 to 0) := (others => '0');
    variable r2246 : std_logic_vector(0 to 0) := (others => '0');
    variable r2245 : std_logic_vector(0 to 0) := (others => '0');
    variable r2244 : std_logic_vector(0 to 0) := (others => '0');
    variable r2243 : std_logic_vector(0 to 0) := (others => '0');
    variable r2242 : std_logic_vector(0 to 0) := (others => '0');
    variable r2241 : std_logic_vector(0 to 0) := (others => '0');
    variable r2240 : std_logic_vector(0 to 0) := (others => '0');
    variable r2239 : std_logic_vector(0 to 0) := (others => '0');
    variable r2238 : std_logic_vector(0 to 0) := (others => '0');
    variable r2237 : std_logic_vector(0 to 0) := (others => '0');
    variable r2236 : std_logic_vector(0 to 0) := (others => '0');
    variable r2235 : std_logic_vector(0 to 0) := (others => '0');
    variable r2234 : std_logic_vector(0 to 0) := (others => '0');
    variable r2233 : std_logic_vector(0 to 0) := (others => '0');
    variable r2232 : std_logic_vector(0 to 0) := (others => '0');
    variable r2231 : std_logic_vector(0 to 0) := (others => '0');
    variable r2230 : std_logic_vector(0 to 0) := (others => '0');
    variable r2229 : std_logic_vector(0 to 0) := (others => '0');
    variable r2228 : std_logic_vector(0 to 0) := (others => '0');
    variable r2227 : std_logic_vector(0 to 0) := (others => '0');
    variable r2226 : std_logic_vector(0 to 0) := (others => '0');
    variable r2225 : std_logic_vector(0 to 0) := (others => '0');
    variable r2224 : std_logic_vector(0 to 0) := (others => '0');
    variable r2223 : std_logic_vector(0 to 0) := (others => '0');
    variable r2222 : std_logic_vector(0 to 0) := (others => '0');
    variable b2221 : boolean := false;
    variable r2220 : std_logic_vector(0 to 31) := (others => '0');
  begin
    b2221 := true;
    r2222 := r2218(0 to 0);
    r2223 := r2218(1 to 1);
    r2224 := r2218(2 to 2);
    r2225 := r2218(3 to 3);
    r2226 := r2218(4 to 4);
    r2227 := r2218(5 to 5);
    r2228 := r2218(6 to 6);
    r2229 := r2218(7 to 7);
    r2230 := r2218(8 to 8);
    r2231 := r2218(9 to 9);
    r2232 := r2218(10 to 10);
    r2233 := r2218(11 to 11);
    r2234 := r2218(12 to 12);
    r2235 := r2218(13 to 13);
    r2236 := r2218(14 to 14);
    r2237 := r2218(15 to 15);
    r2238 := r2218(16 to 16);
    r2239 := r2218(17 to 17);
    r2240 := r2218(18 to 18);
    r2241 := r2218(19 to 19);
    r2242 := r2218(20 to 20);
    r2243 := r2218(21 to 21);
    r2244 := r2218(22 to 22);
    r2245 := r2218(23 to 23);
    r2246 := r2218(24 to 24);
    r2247 := r2218(25 to 25);
    r2248 := r2218(26 to 26);
    r2249 := r2218(27 to 27);
    r2250 := r2218(28 to 28);
    r2251 := r2218(29 to 29);
    r2252 := r2218(30 to 30);
    r2253 := r2218(31 to 31);
    b2254 := true;
    b2255 := true;
    b2256 := true;
    b2257 := true;
    b2258 := true;
    b2259 := true;
    b2260 := true;
    b2261 := true;
    b2262 := true;
    b2263 := true;
    b2264 := true;
    b2265 := true;
    b2266 := true;
    b2267 := true;
    b2268 := true;
    b2269 := true;
    b2270 := true;
    b2271 := true;
    b2272 := true;
    b2273 := true;
    b2274 := true;
    b2275 := true;
    b2276 := true;
    b2277 := true;
    b2278 := true;
    b2279 := true;
    b2280 := true;
    b2281 := true;
    b2282 := true;
    b2283 := true;
    b2284 := true;
    b2285 := true;
    b2286 := (b2254 AND (b2255 AND (b2256 AND (b2257 AND (b2258 AND (b2259 AND (b2260 AND (b2261 AND (b2262 AND (b2263 AND (b2264 AND (b2265 AND (b2266 AND (b2267 AND (b2268 AND (b2269 AND (b2270 AND (b2271 AND (b2272 AND (b2273 AND (b2274 AND (b2275 AND (b2276 AND (b2277 AND (b2278 AND (b2279 AND (b2280 AND (b2281 AND (b2282 AND (b2283 AND (b2284 AND b2285)))))))))))))))))))))))))))))));
    if b2286 then
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      r2288 := (r2241 & r2242 & r2243 & r2244 & r2245 & r2246 & r2247 & r2248 & r2249 & r2250 & r2251 & r2252 & r2253 & r2222 & r2223 & r2224 & r2225 & r2226 & r2227 & r2228 & r2229 & r2230 & r2231 & r2232 & r2233 & r2234 & r2235 & r2236 & r2237 & r2238 & r2239 & r2240);
      r2220 := r2288;
    end if;
    return r2220;
  end rewire_rot13_2217;
  function rewire_rot9_2142(r2143 : std_logic_vector) return std_logic_vector
  is
    variable r2213 : std_logic_vector(0 to 31) := (others => '0');
    variable EMPTY : std_logic_vector(0 to -1) := (others => '0');
    variable b2211 : boolean := false;
    variable b2210 : boolean := false;
    variable b2209 : boolean := false;
    variable b2208 : boolean := false;
    variable b2207 : boolean := false;
    variable b2206 : boolean := false;
    variable b2205 : boolean := false;
    variable b2204 : boolean := false;
    variable b2203 : boolean := false;
    variable b2202 : boolean := false;
    variable b2201 : boolean := false;
    variable b2200 : boolean := false;
    variable b2199 : boolean := false;
    variable b2198 : boolean := false;
    variable b2197 : boolean := false;
    variable b2196 : boolean := false;
    variable b2195 : boolean := false;
    variable b2194 : boolean := false;
    variable b2193 : boolean := false;
    variable b2192 : boolean := false;
    variable b2191 : boolean := false;
    variable b2190 : boolean := false;
    variable b2189 : boolean := false;
    variable b2188 : boolean := false;
    variable b2187 : boolean := false;
    variable b2186 : boolean := false;
    variable b2185 : boolean := false;
    variable b2184 : boolean := false;
    variable b2183 : boolean := false;
    variable b2182 : boolean := false;
    variable b2181 : boolean := false;
    variable b2180 : boolean := false;
    variable b2179 : boolean := false;
    variable r2178 : std_logic_vector(0 to 0) := (others => '0');
    variable r2177 : std_logic_vector(0 to 0) := (others => '0');
    variable r2176 : std_logic_vector(0 to 0) := (others => '0');
    variable r2175 : std_logic_vector(0 to 0) := (others => '0');
    variable r2174 : std_logic_vector(0 to 0) := (others => '0');
    variable r2173 : std_logic_vector(0 to 0) := (others => '0');
    variable r2172 : std_logic_vector(0 to 0) := (others => '0');
    variable r2171 : std_logic_vector(0 to 0) := (others => '0');
    variable r2170 : std_logic_vector(0 to 0) := (others => '0');
    variable r2169 : std_logic_vector(0 to 0) := (others => '0');
    variable r2168 : std_logic_vector(0 to 0) := (others => '0');
    variable r2167 : std_logic_vector(0 to 0) := (others => '0');
    variable r2166 : std_logic_vector(0 to 0) := (others => '0');
    variable r2165 : std_logic_vector(0 to 0) := (others => '0');
    variable r2164 : std_logic_vector(0 to 0) := (others => '0');
    variable r2163 : std_logic_vector(0 to 0) := (others => '0');
    variable r2162 : std_logic_vector(0 to 0) := (others => '0');
    variable r2161 : std_logic_vector(0 to 0) := (others => '0');
    variable r2160 : std_logic_vector(0 to 0) := (others => '0');
    variable r2159 : std_logic_vector(0 to 0) := (others => '0');
    variable r2158 : std_logic_vector(0 to 0) := (others => '0');
    variable r2157 : std_logic_vector(0 to 0) := (others => '0');
    variable r2156 : std_logic_vector(0 to 0) := (others => '0');
    variable r2155 : std_logic_vector(0 to 0) := (others => '0');
    variable r2154 : std_logic_vector(0 to 0) := (others => '0');
    variable r2153 : std_logic_vector(0 to 0) := (others => '0');
    variable r2152 : std_logic_vector(0 to 0) := (others => '0');
    variable r2151 : std_logic_vector(0 to 0) := (others => '0');
    variable r2150 : std_logic_vector(0 to 0) := (others => '0');
    variable r2149 : std_logic_vector(0 to 0) := (others => '0');
    variable r2148 : std_logic_vector(0 to 0) := (others => '0');
    variable r2147 : std_logic_vector(0 to 0) := (others => '0');
    variable b2146 : boolean := false;
    variable r2145 : std_logic_vector(0 to 31) := (others => '0');
  begin
    b2146 := true;
    r2147 := r2143(0 to 0);
    r2148 := r2143(1 to 1);
    r2149 := r2143(2 to 2);
    r2150 := r2143(3 to 3);
    r2151 := r2143(4 to 4);
    r2152 := r2143(5 to 5);
    r2153 := r2143(6 to 6);
    r2154 := r2143(7 to 7);
    r2155 := r2143(8 to 8);
    r2156 := r2143(9 to 9);
    r2157 := r2143(10 to 10);
    r2158 := r2143(11 to 11);
    r2159 := r2143(12 to 12);
    r2160 := r2143(13 to 13);
    r2161 := r2143(14 to 14);
    r2162 := r2143(15 to 15);
    r2163 := r2143(16 to 16);
    r2164 := r2143(17 to 17);
    r2165 := r2143(18 to 18);
    r2166 := r2143(19 to 19);
    r2167 := r2143(20 to 20);
    r2168 := r2143(21 to 21);
    r2169 := r2143(22 to 22);
    r2170 := r2143(23 to 23);
    r2171 := r2143(24 to 24);
    r2172 := r2143(25 to 25);
    r2173 := r2143(26 to 26);
    r2174 := r2143(27 to 27);
    r2175 := r2143(28 to 28);
    r2176 := r2143(29 to 29);
    r2177 := r2143(30 to 30);
    r2178 := r2143(31 to 31);
    b2179 := true;
    b2180 := true;
    b2181 := true;
    b2182 := true;
    b2183 := true;
    b2184 := true;
    b2185 := true;
    b2186 := true;
    b2187 := true;
    b2188 := true;
    b2189 := true;
    b2190 := true;
    b2191 := true;
    b2192 := true;
    b2193 := true;
    b2194 := true;
    b2195 := true;
    b2196 := true;
    b2197 := true;
    b2198 := true;
    b2199 := true;
    b2200 := true;
    b2201 := true;
    b2202 := true;
    b2203 := true;
    b2204 := true;
    b2205 := true;
    b2206 := true;
    b2207 := true;
    b2208 := true;
    b2209 := true;
    b2210 := true;
    b2211 := (b2179 AND (b2180 AND (b2181 AND (b2182 AND (b2183 AND (b2184 AND (b2185 AND (b2186 AND (b2187 AND (b2188 AND (b2189 AND (b2190 AND (b2191 AND (b2192 AND (b2193 AND (b2194 AND (b2195 AND (b2196 AND (b2197 AND (b2198 AND (b2199 AND (b2200 AND (b2201 AND (b2202 AND (b2203 AND (b2204 AND (b2205 AND (b2206 AND (b2207 AND (b2208 AND (b2209 AND b2210)))))))))))))))))))))))))))))));
    if b2211 then
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      r2213 := (r2170 & r2171 & r2172 & r2173 & r2174 & r2175 & r2176 & r2177 & r2178 & r2147 & r2148 & r2149 & r2150 & r2151 & r2152 & r2153 & r2154 & r2155 & r2156 & r2157 & r2158 & r2159 & r2160 & r2161 & r2162 & r2163 & r2164 & r2165 & r2166 & r2167 & r2168 & r2169);
      r2145 := r2213;
    end if;
    return r2145;
  end rewire_rot9_2142;
  function rewire_rot7_2067(r2068 : std_logic_vector) return std_logic_vector
  is
    variable r2138 : std_logic_vector(0 to 31) := (others => '0');
    variable EMPTY : std_logic_vector(0 to -1) := (others => '0');
    variable b2136 : boolean := false;
    variable b2135 : boolean := false;
    variable b2134 : boolean := false;
    variable b2133 : boolean := false;
    variable b2132 : boolean := false;
    variable b2131 : boolean := false;
    variable b2130 : boolean := false;
    variable b2129 : boolean := false;
    variable b2128 : boolean := false;
    variable b2127 : boolean := false;
    variable b2126 : boolean := false;
    variable b2125 : boolean := false;
    variable b2124 : boolean := false;
    variable b2123 : boolean := false;
    variable b2122 : boolean := false;
    variable b2121 : boolean := false;
    variable b2120 : boolean := false;
    variable b2119 : boolean := false;
    variable b2118 : boolean := false;
    variable b2117 : boolean := false;
    variable b2116 : boolean := false;
    variable b2115 : boolean := false;
    variable b2114 : boolean := false;
    variable b2113 : boolean := false;
    variable b2112 : boolean := false;
    variable b2111 : boolean := false;
    variable b2110 : boolean := false;
    variable b2109 : boolean := false;
    variable b2108 : boolean := false;
    variable b2107 : boolean := false;
    variable b2106 : boolean := false;
    variable b2105 : boolean := false;
    variable b2104 : boolean := false;
    variable r2103 : std_logic_vector(0 to 0) := (others => '0');
    variable r2102 : std_logic_vector(0 to 0) := (others => '0');
    variable r2101 : std_logic_vector(0 to 0) := (others => '0');
    variable r2100 : std_logic_vector(0 to 0) := (others => '0');
    variable r2099 : std_logic_vector(0 to 0) := (others => '0');
    variable r2098 : std_logic_vector(0 to 0) := (others => '0');
    variable r2097 : std_logic_vector(0 to 0) := (others => '0');
    variable r2096 : std_logic_vector(0 to 0) := (others => '0');
    variable r2095 : std_logic_vector(0 to 0) := (others => '0');
    variable r2094 : std_logic_vector(0 to 0) := (others => '0');
    variable r2093 : std_logic_vector(0 to 0) := (others => '0');
    variable r2092 : std_logic_vector(0 to 0) := (others => '0');
    variable r2091 : std_logic_vector(0 to 0) := (others => '0');
    variable r2090 : std_logic_vector(0 to 0) := (others => '0');
    variable r2089 : std_logic_vector(0 to 0) := (others => '0');
    variable r2088 : std_logic_vector(0 to 0) := (others => '0');
    variable r2087 : std_logic_vector(0 to 0) := (others => '0');
    variable r2086 : std_logic_vector(0 to 0) := (others => '0');
    variable r2085 : std_logic_vector(0 to 0) := (others => '0');
    variable r2084 : std_logic_vector(0 to 0) := (others => '0');
    variable r2083 : std_logic_vector(0 to 0) := (others => '0');
    variable r2082 : std_logic_vector(0 to 0) := (others => '0');
    variable r2081 : std_logic_vector(0 to 0) := (others => '0');
    variable r2080 : std_logic_vector(0 to 0) := (others => '0');
    variable r2079 : std_logic_vector(0 to 0) := (others => '0');
    variable r2078 : std_logic_vector(0 to 0) := (others => '0');
    variable r2077 : std_logic_vector(0 to 0) := (others => '0');
    variable r2076 : std_logic_vector(0 to 0) := (others => '0');
    variable r2075 : std_logic_vector(0 to 0) := (others => '0');
    variable r2074 : std_logic_vector(0 to 0) := (others => '0');
    variable r2073 : std_logic_vector(0 to 0) := (others => '0');
    variable r2072 : std_logic_vector(0 to 0) := (others => '0');
    variable b2071 : boolean := false;
    variable r2070 : std_logic_vector(0 to 31) := (others => '0');
  begin
    b2071 := true;
    r2072 := r2068(0 to 0);
    r2073 := r2068(1 to 1);
    r2074 := r2068(2 to 2);
    r2075 := r2068(3 to 3);
    r2076 := r2068(4 to 4);
    r2077 := r2068(5 to 5);
    r2078 := r2068(6 to 6);
    r2079 := r2068(7 to 7);
    r2080 := r2068(8 to 8);
    r2081 := r2068(9 to 9);
    r2082 := r2068(10 to 10);
    r2083 := r2068(11 to 11);
    r2084 := r2068(12 to 12);
    r2085 := r2068(13 to 13);
    r2086 := r2068(14 to 14);
    r2087 := r2068(15 to 15);
    r2088 := r2068(16 to 16);
    r2089 := r2068(17 to 17);
    r2090 := r2068(18 to 18);
    r2091 := r2068(19 to 19);
    r2092 := r2068(20 to 20);
    r2093 := r2068(21 to 21);
    r2094 := r2068(22 to 22);
    r2095 := r2068(23 to 23);
    r2096 := r2068(24 to 24);
    r2097 := r2068(25 to 25);
    r2098 := r2068(26 to 26);
    r2099 := r2068(27 to 27);
    r2100 := r2068(28 to 28);
    r2101 := r2068(29 to 29);
    r2102 := r2068(30 to 30);
    r2103 := r2068(31 to 31);
    b2104 := true;
    b2105 := true;
    b2106 := true;
    b2107 := true;
    b2108 := true;
    b2109 := true;
    b2110 := true;
    b2111 := true;
    b2112 := true;
    b2113 := true;
    b2114 := true;
    b2115 := true;
    b2116 := true;
    b2117 := true;
    b2118 := true;
    b2119 := true;
    b2120 := true;
    b2121 := true;
    b2122 := true;
    b2123 := true;
    b2124 := true;
    b2125 := true;
    b2126 := true;
    b2127 := true;
    b2128 := true;
    b2129 := true;
    b2130 := true;
    b2131 := true;
    b2132 := true;
    b2133 := true;
    b2134 := true;
    b2135 := true;
    b2136 := (b2104 AND (b2105 AND (b2106 AND (b2107 AND (b2108 AND (b2109 AND (b2110 AND (b2111 AND (b2112 AND (b2113 AND (b2114 AND (b2115 AND (b2116 AND (b2117 AND (b2118 AND (b2119 AND (b2120 AND (b2121 AND (b2122 AND (b2123 AND (b2124 AND (b2125 AND (b2126 AND (b2127 AND (b2128 AND (b2129 AND (b2130 AND (b2131 AND (b2132 AND (b2133 AND (b2134 AND b2135)))))))))))))))))))))))))))))));
    if b2136 then
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      r2138 := (r2097 & r2098 & r2099 & r2100 & r2101 & r2102 & r2103 & r2072 & r2073 & r2074 & r2075 & r2076 & r2077 & r2078 & r2079 & r2080 & r2081 & r2082 & r2083 & r2084 & r2085 & r2086 & r2087 & r2088 & r2089 & r2090 & r2091 & r2092 & r2093 & r2094 & r2095 & r2096);
      r2070 := r2138;
    end if;
    return r2070;
  end rewire_rot7_2067;
  function rewire_expwords_1657(r1658 : std_logic_vector) return std_logic_vector
  is
    variable r1973 : std_logic_vector(0 to 511) := (others => '0');
    variable b1971 : boolean := false;
    variable b1970 : boolean := false;
    variable b1969 : boolean := false;
    variable b1968 : boolean := false;
    variable b1967 : boolean := false;
    variable b1966 : boolean := false;
    variable r1965 : std_logic_vector(0 to 7) := (others => '0');
    variable r1964 : std_logic_vector(0 to 7) := (others => '0');
    variable r1963 : std_logic_vector(0 to 7) := (others => '0');
    variable r1962 : std_logic_vector(0 to 7) := (others => '0');
    variable b1961 : boolean := false;
    variable b1960 : boolean := false;
    variable b1959 : boolean := false;
    variable b1958 : boolean := false;
    variable b1957 : boolean := false;
    variable b1956 : boolean := false;
    variable r1955 : std_logic_vector(0 to 7) := (others => '0');
    variable r1954 : std_logic_vector(0 to 7) := (others => '0');
    variable r1953 : std_logic_vector(0 to 7) := (others => '0');
    variable r1952 : std_logic_vector(0 to 7) := (others => '0');
    variable b1951 : boolean := false;
    variable b1950 : boolean := false;
    variable b1949 : boolean := false;
    variable b1948 : boolean := false;
    variable b1947 : boolean := false;
    variable b1946 : boolean := false;
    variable r1945 : std_logic_vector(0 to 7) := (others => '0');
    variable r1944 : std_logic_vector(0 to 7) := (others => '0');
    variable r1943 : std_logic_vector(0 to 7) := (others => '0');
    variable r1942 : std_logic_vector(0 to 7) := (others => '0');
    variable b1941 : boolean := false;
    variable b1940 : boolean := false;
    variable b1939 : boolean := false;
    variable b1938 : boolean := false;
    variable b1937 : boolean := false;
    variable b1936 : boolean := false;
    variable r1935 : std_logic_vector(0 to 7) := (others => '0');
    variable r1934 : std_logic_vector(0 to 7) := (others => '0');
    variable r1933 : std_logic_vector(0 to 7) := (others => '0');
    variable r1932 : std_logic_vector(0 to 7) := (others => '0');
    variable b1931 : boolean := false;
    variable b1930 : boolean := false;
    variable b1929 : boolean := false;
    variable b1928 : boolean := false;
    variable b1927 : boolean := false;
    variable b1926 : boolean := false;
    variable r1925 : std_logic_vector(0 to 7) := (others => '0');
    variable r1924 : std_logic_vector(0 to 7) := (others => '0');
    variable r1923 : std_logic_vector(0 to 7) := (others => '0');
    variable r1922 : std_logic_vector(0 to 7) := (others => '0');
    variable b1921 : boolean := false;
    variable b1920 : boolean := false;
    variable b1919 : boolean := false;
    variable b1918 : boolean := false;
    variable b1917 : boolean := false;
    variable b1916 : boolean := false;
    variable r1915 : std_logic_vector(0 to 7) := (others => '0');
    variable r1914 : std_logic_vector(0 to 7) := (others => '0');
    variable r1913 : std_logic_vector(0 to 7) := (others => '0');
    variable r1912 : std_logic_vector(0 to 7) := (others => '0');
    variable b1911 : boolean := false;
    variable b1910 : boolean := false;
    variable b1909 : boolean := false;
    variable b1908 : boolean := false;
    variable b1907 : boolean := false;
    variable b1906 : boolean := false;
    variable r1905 : std_logic_vector(0 to 7) := (others => '0');
    variable r1904 : std_logic_vector(0 to 7) := (others => '0');
    variable r1903 : std_logic_vector(0 to 7) := (others => '0');
    variable r1902 : std_logic_vector(0 to 7) := (others => '0');
    variable b1901 : boolean := false;
    variable b1900 : boolean := false;
    variable b1899 : boolean := false;
    variable b1898 : boolean := false;
    variable b1897 : boolean := false;
    variable b1896 : boolean := false;
    variable r1895 : std_logic_vector(0 to 7) := (others => '0');
    variable r1894 : std_logic_vector(0 to 7) := (others => '0');
    variable r1893 : std_logic_vector(0 to 7) := (others => '0');
    variable r1892 : std_logic_vector(0 to 7) := (others => '0');
    variable b1891 : boolean := false;
    variable b1890 : boolean := false;
    variable b1889 : boolean := false;
    variable b1888 : boolean := false;
    variable b1887 : boolean := false;
    variable b1886 : boolean := false;
    variable r1885 : std_logic_vector(0 to 7) := (others => '0');
    variable r1884 : std_logic_vector(0 to 7) := (others => '0');
    variable r1883 : std_logic_vector(0 to 7) := (others => '0');
    variable r1882 : std_logic_vector(0 to 7) := (others => '0');
    variable b1881 : boolean := false;
    variable b1880 : boolean := false;
    variable b1879 : boolean := false;
    variable b1878 : boolean := false;
    variable b1877 : boolean := false;
    variable b1876 : boolean := false;
    variable r1875 : std_logic_vector(0 to 7) := (others => '0');
    variable r1874 : std_logic_vector(0 to 7) := (others => '0');
    variable r1873 : std_logic_vector(0 to 7) := (others => '0');
    variable r1872 : std_logic_vector(0 to 7) := (others => '0');
    variable b1871 : boolean := false;
    variable b1870 : boolean := false;
    variable b1869 : boolean := false;
    variable b1868 : boolean := false;
    variable b1867 : boolean := false;
    variable b1866 : boolean := false;
    variable r1865 : std_logic_vector(0 to 7) := (others => '0');
    variable r1864 : std_logic_vector(0 to 7) := (others => '0');
    variable r1863 : std_logic_vector(0 to 7) := (others => '0');
    variable r1862 : std_logic_vector(0 to 7) := (others => '0');
    variable b1861 : boolean := false;
    variable b1860 : boolean := false;
    variable b1859 : boolean := false;
    variable b1858 : boolean := false;
    variable b1857 : boolean := false;
    variable b1856 : boolean := false;
    variable r1855 : std_logic_vector(0 to 7) := (others => '0');
    variable r1854 : std_logic_vector(0 to 7) := (others => '0');
    variable r1853 : std_logic_vector(0 to 7) := (others => '0');
    variable r1852 : std_logic_vector(0 to 7) := (others => '0');
    variable b1851 : boolean := false;
    variable b1850 : boolean := false;
    variable b1849 : boolean := false;
    variable b1848 : boolean := false;
    variable b1847 : boolean := false;
    variable b1846 : boolean := false;
    variable r1845 : std_logic_vector(0 to 7) := (others => '0');
    variable r1844 : std_logic_vector(0 to 7) := (others => '0');
    variable r1843 : std_logic_vector(0 to 7) := (others => '0');
    variable r1842 : std_logic_vector(0 to 7) := (others => '0');
    variable b1841 : boolean := false;
    variable b1840 : boolean := false;
    variable b1839 : boolean := false;
    variable b1838 : boolean := false;
    variable b1837 : boolean := false;
    variable b1836 : boolean := false;
    variable r1835 : std_logic_vector(0 to 7) := (others => '0');
    variable r1834 : std_logic_vector(0 to 7) := (others => '0');
    variable r1833 : std_logic_vector(0 to 7) := (others => '0');
    variable r1832 : std_logic_vector(0 to 7) := (others => '0');
    variable b1831 : boolean := false;
    variable b1830 : boolean := false;
    variable b1829 : boolean := false;
    variable b1828 : boolean := false;
    variable b1827 : boolean := false;
    variable b1826 : boolean := false;
    variable r1825 : std_logic_vector(0 to 7) := (others => '0');
    variable r1824 : std_logic_vector(0 to 7) := (others => '0');
    variable r1823 : std_logic_vector(0 to 7) := (others => '0');
    variable r1822 : std_logic_vector(0 to 7) := (others => '0');
    variable b1821 : boolean := false;
    variable b1820 : boolean := false;
    variable b1819 : boolean := false;
    variable b1818 : boolean := false;
    variable b1817 : boolean := false;
    variable b1816 : boolean := false;
    variable r1815 : std_logic_vector(0 to 7) := (others => '0');
    variable r1814 : std_logic_vector(0 to 7) := (others => '0');
    variable r1813 : std_logic_vector(0 to 7) := (others => '0');
    variable r1812 : std_logic_vector(0 to 7) := (others => '0');
    variable b1811 : boolean := false;
    variable r1810 : std_logic_vector(0 to 31) := (others => '0');
    variable r1809 : std_logic_vector(0 to 31) := (others => '0');
    variable r1808 : std_logic_vector(0 to 31) := (others => '0');
    variable r1807 : std_logic_vector(0 to 31) := (others => '0');
    variable r1806 : std_logic_vector(0 to 31) := (others => '0');
    variable r1805 : std_logic_vector(0 to 31) := (others => '0');
    variable r1804 : std_logic_vector(0 to 31) := (others => '0');
    variable r1803 : std_logic_vector(0 to 31) := (others => '0');
    variable r1802 : std_logic_vector(0 to 31) := (others => '0');
    variable r1801 : std_logic_vector(0 to 31) := (others => '0');
    variable r1800 : std_logic_vector(0 to 31) := (others => '0');
    variable r1799 : std_logic_vector(0 to 31) := (others => '0');
    variable r1798 : std_logic_vector(0 to 31) := (others => '0');
    variable r1797 : std_logic_vector(0 to 31) := (others => '0');
    variable r1796 : std_logic_vector(0 to 31) := (others => '0');
    variable r1795 : std_logic_vector(0 to 31) := (others => '0');
    variable b1794 : boolean := false;
    variable r1793 : std_logic_vector(0 to 511) := (others => '0');
    variable r1792 : std_logic_vector(0 to 511) := (others => '0');
    variable EMPTY : std_logic_vector(0 to -1) := (others => '0');
    variable r1790 : std_logic_vector(0 to 31) := (others => '0');
    variable r1789 : std_logic_vector(0 to 31) := (others => '0');
    variable r1788 : std_logic_vector(0 to 31) := (others => '0');
    variable r1787 : std_logic_vector(0 to 31) := (others => '0');
    variable r1786 : std_logic_vector(0 to 31) := (others => '0');
    variable r1785 : std_logic_vector(0 to 31) := (others => '0');
    variable r1784 : std_logic_vector(0 to 31) := (others => '0');
    variable r1783 : std_logic_vector(0 to 31) := (others => '0');
    variable r1782 : std_logic_vector(0 to 31) := (others => '0');
    variable r1781 : std_logic_vector(0 to 31) := (others => '0');
    variable r1780 : std_logic_vector(0 to 31) := (others => '0');
    variable r1779 : std_logic_vector(0 to 31) := (others => '0');
    variable r1778 : std_logic_vector(0 to 31) := (others => '0');
    variable r1777 : std_logic_vector(0 to 31) := (others => '0');
    variable r1776 : std_logic_vector(0 to 31) := (others => '0');
    variable r1775 : std_logic_vector(0 to 31) := (others => '0');
    variable r1697 : std_logic_vector(0 to 31) := (others => '0');
    variable r1696 : std_logic_vector(0 to 31) := (others => '0');
    variable b1694 : boolean := false;
    variable b1693 : boolean := false;
    variable b1692 : boolean := false;
    variable b1691 : boolean := false;
    variable b1690 : boolean := false;
    variable b1689 : boolean := false;
    variable b1688 : boolean := false;
    variable b1687 : boolean := false;
    variable b1686 : boolean := false;
    variable b1685 : boolean := false;
    variable b1684 : boolean := false;
    variable b1683 : boolean := false;
    variable b1682 : boolean := false;
    variable b1681 : boolean := false;
    variable b1680 : boolean := false;
    variable b1679 : boolean := false;
    variable b1678 : boolean := false;
    variable r1677 : std_logic_vector(0 to 31) := (others => '0');
    variable r1676 : std_logic_vector(0 to 31) := (others => '0');
    variable r1675 : std_logic_vector(0 to 31) := (others => '0');
    variable r1674 : std_logic_vector(0 to 31) := (others => '0');
    variable r1673 : std_logic_vector(0 to 31) := (others => '0');
    variable r1672 : std_logic_vector(0 to 31) := (others => '0');
    variable r1671 : std_logic_vector(0 to 31) := (others => '0');
    variable r1670 : std_logic_vector(0 to 31) := (others => '0');
    variable r1669 : std_logic_vector(0 to 31) := (others => '0');
    variable r1668 : std_logic_vector(0 to 31) := (others => '0');
    variable r1667 : std_logic_vector(0 to 31) := (others => '0');
    variable r1666 : std_logic_vector(0 to 31) := (others => '0');
    variable r1665 : std_logic_vector(0 to 31) := (others => '0');
    variable r1664 : std_logic_vector(0 to 31) := (others => '0');
    variable r1663 : std_logic_vector(0 to 31) := (others => '0');
    variable r1662 : std_logic_vector(0 to 31) := (others => '0');
    variable b1661 : boolean := false;
    variable r1660 : std_logic_vector(0 to 511) := (others => '0');
  begin
    b1661 := true;
    r1662 := r1658(0 to 31);
    r1663 := r1658(32 to 63);
    r1664 := r1658(64 to 95);
    r1665 := r1658(96 to 127);
    r1666 := r1658(128 to 159);
    r1667 := r1658(160 to 191);
    r1668 := r1658(192 to 223);
    r1669 := r1658(224 to 255);
    r1670 := r1658(256 to 287);
    r1671 := r1658(288 to 319);
    r1672 := r1658(320 to 351);
    r1673 := r1658(352 to 383);
    r1674 := r1658(384 to 415);
    r1675 := r1658(416 to 447);
    r1676 := r1658(448 to 479);
    r1677 := r1658(480 to 511);
    b1678 := true;
    b1679 := true;
    b1680 := true;
    b1681 := true;
    b1682 := true;
    b1683 := true;
    b1684 := true;
    b1685 := true;
    b1686 := true;
    b1687 := true;
    b1688 := true;
    b1689 := true;
    b1690 := true;
    b1691 := true;
    b1692 := true;
    b1693 := true;
    b1694 := (b1678 AND (b1679 AND (b1680 AND (b1681 AND (b1682 AND (b1683 AND (b1684 AND (b1685 AND (b1686 AND (b1687 AND (b1688 AND (b1689 AND (b1690 AND (b1691 AND (b1692 AND b1693)))))))))))))));
    if b1694 then
      null;
      r1775 := rewire_littleendianp_1695(r1662);
      null;
      r1776 := rewire_littleendianp_1695(r1663);
      null;
      r1777 := rewire_littleendianp_1695(r1664);
      null;
      r1778 := rewire_littleendianp_1695(r1665);
      null;
      r1779 := rewire_littleendianp_1695(r1666);
      null;
      r1780 := rewire_littleendianp_1695(r1667);
      null;
      r1781 := rewire_littleendianp_1695(r1668);
      null;
      r1782 := rewire_littleendianp_1695(r1669);
      null;
      r1783 := rewire_littleendianp_1695(r1670);
      null;
      r1784 := rewire_littleendianp_1695(r1671);
      null;
      r1785 := rewire_littleendianp_1695(r1672);
      null;
      r1786 := rewire_littleendianp_1695(r1673);
      null;
      r1787 := rewire_littleendianp_1695(r1674);
      null;
      r1788 := rewire_littleendianp_1695(r1675);
      null;
      r1789 := rewire_littleendianp_1695(r1676);
      null;
      r1790 := rewire_littleendianp_1695(r1677);
      b1794 := true;
      r1795 := r1792(0 to 31);
      r1796 := r1792(32 to 63);
      r1797 := r1792(64 to 95);
      r1798 := r1792(96 to 127);
      r1799 := r1792(128 to 159);
      r1800 := r1792(160 to 191);
      r1801 := r1792(192 to 223);
      r1802 := r1792(224 to 255);
      r1803 := r1792(256 to 287);
      r1804 := r1792(288 to 319);
      r1805 := r1792(320 to 351);
      r1806 := r1792(352 to 383);
      r1807 := r1792(384 to 415);
      r1808 := r1792(416 to 447);
      r1809 := r1792(448 to 479);
      r1810 := r1792(480 to 511);
      b1811 := true;
      r1812 := r1795(0 to 7);
      r1813 := r1795(8 to 15);
      r1814 := r1795(16 to 23);
      r1815 := r1795(24 to 31);
      b1816 := true;
      b1817 := true;
      b1818 := true;
      b1819 := true;
      b1820 := (b1816 AND (b1817 AND (b1818 AND b1819)));
      b1821 := true;
      r1822 := r1796(0 to 7);
      r1823 := r1796(8 to 15);
      r1824 := r1796(16 to 23);
      r1825 := r1796(24 to 31);
      b1826 := true;
      b1827 := true;
      b1828 := true;
      b1829 := true;
      b1830 := (b1826 AND (b1827 AND (b1828 AND b1829)));
      b1831 := true;
      r1832 := r1797(0 to 7);
      r1833 := r1797(8 to 15);
      r1834 := r1797(16 to 23);
      r1835 := r1797(24 to 31);
      b1836 := true;
      b1837 := true;
      b1838 := true;
      b1839 := true;
      b1840 := (b1836 AND (b1837 AND (b1838 AND b1839)));
      b1841 := true;
      r1842 := r1798(0 to 7);
      r1843 := r1798(8 to 15);
      r1844 := r1798(16 to 23);
      r1845 := r1798(24 to 31);
      b1846 := true;
      b1847 := true;
      b1848 := true;
      b1849 := true;
      b1850 := (b1846 AND (b1847 AND (b1848 AND b1849)));
      b1851 := true;
      r1852 := r1799(0 to 7);
      r1853 := r1799(8 to 15);
      r1854 := r1799(16 to 23);
      r1855 := r1799(24 to 31);
      b1856 := true;
      b1857 := true;
      b1858 := true;
      b1859 := true;
      b1860 := (b1856 AND (b1857 AND (b1858 AND b1859)));
      b1861 := true;
      r1862 := r1800(0 to 7);
      r1863 := r1800(8 to 15);
      r1864 := r1800(16 to 23);
      r1865 := r1800(24 to 31);
      b1866 := true;
      b1867 := true;
      b1868 := true;
      b1869 := true;
      b1870 := (b1866 AND (b1867 AND (b1868 AND b1869)));
      b1871 := true;
      r1872 := r1801(0 to 7);
      r1873 := r1801(8 to 15);
      r1874 := r1801(16 to 23);
      r1875 := r1801(24 to 31);
      b1876 := true;
      b1877 := true;
      b1878 := true;
      b1879 := true;
      b1880 := (b1876 AND (b1877 AND (b1878 AND b1879)));
      b1881 := true;
      r1882 := r1802(0 to 7);
      r1883 := r1802(8 to 15);
      r1884 := r1802(16 to 23);
      r1885 := r1802(24 to 31);
      b1886 := true;
      b1887 := true;
      b1888 := true;
      b1889 := true;
      b1890 := (b1886 AND (b1887 AND (b1888 AND b1889)));
      b1891 := true;
      r1892 := r1803(0 to 7);
      r1893 := r1803(8 to 15);
      r1894 := r1803(16 to 23);
      r1895 := r1803(24 to 31);
      b1896 := true;
      b1897 := true;
      b1898 := true;
      b1899 := true;
      b1900 := (b1896 AND (b1897 AND (b1898 AND b1899)));
      b1901 := true;
      r1902 := r1804(0 to 7);
      r1903 := r1804(8 to 15);
      r1904 := r1804(16 to 23);
      r1905 := r1804(24 to 31);
      b1906 := true;
      b1907 := true;
      b1908 := true;
      b1909 := true;
      b1910 := (b1906 AND (b1907 AND (b1908 AND b1909)));
      b1911 := true;
      r1912 := r1805(0 to 7);
      r1913 := r1805(8 to 15);
      r1914 := r1805(16 to 23);
      r1915 := r1805(24 to 31);
      b1916 := true;
      b1917 := true;
      b1918 := true;
      b1919 := true;
      b1920 := (b1916 AND (b1917 AND (b1918 AND b1919)));
      b1921 := true;
      r1922 := r1806(0 to 7);
      r1923 := r1806(8 to 15);
      r1924 := r1806(16 to 23);
      r1925 := r1806(24 to 31);
      b1926 := true;
      b1927 := true;
      b1928 := true;
      b1929 := true;
      b1930 := (b1926 AND (b1927 AND (b1928 AND b1929)));
      b1931 := true;
      r1932 := r1807(0 to 7);
      r1933 := r1807(8 to 15);
      r1934 := r1807(16 to 23);
      r1935 := r1807(24 to 31);
      b1936 := true;
      b1937 := true;
      b1938 := true;
      b1939 := true;
      b1940 := (b1936 AND (b1937 AND (b1938 AND b1939)));
      b1941 := true;
      r1942 := r1808(0 to 7);
      r1943 := r1808(8 to 15);
      r1944 := r1808(16 to 23);
      r1945 := r1808(24 to 31);
      b1946 := true;
      b1947 := true;
      b1948 := true;
      b1949 := true;
      b1950 := (b1946 AND (b1947 AND (b1948 AND b1949)));
      b1951 := true;
      r1952 := r1809(0 to 7);
      r1953 := r1809(8 to 15);
      r1954 := r1809(16 to 23);
      r1955 := r1809(24 to 31);
      b1956 := true;
      b1957 := true;
      b1958 := true;
      b1959 := true;
      b1960 := (b1956 AND (b1957 AND (b1958 AND b1959)));
      b1961 := true;
      r1962 := r1810(0 to 7);
      r1963 := r1810(8 to 15);
      r1964 := r1810(16 to 23);
      r1965 := r1810(24 to 31);
      b1966 := true;
      b1967 := true;
      b1968 := true;
      b1969 := true;
      b1970 := (b1966 AND (b1967 AND (b1968 AND b1969)));
      b1971 := (b1820 AND (b1830 AND (b1840 AND (b1850 AND (b1860 AND (b1870 AND (b1880 AND (b1890 AND (b1900 AND (b1910 AND (b1920 AND (b1930 AND (b1940 AND (b1950 AND (b1960 AND b1970)))))))))))))));
      if b1971 then
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        r1973 := (r1812 & r1813 & r1814 & r1815 & r1822 & r1823 & r1824 & r1825 & r1832 & r1833 & r1834 & r1835 & r1842 & r1843 & r1844 & r1845 & r1852 & r1853 & r1854 & r1855 & r1862 & r1863 & r1864 & r1865 & r1872 & r1873 & r1874 & r1875 & r1882 & r1883 & r1884 & r1885 & r1892 & r1893 & r1894 & r1895 & r1902 & r1903 & r1904 & r1905 & r1912 & r1913 & r1914 & r1915 & r1922 & r1923 & r1924 & r1925 & r1932 & r1933 & r1934 & r1935 & r1942 & r1943 & r1944 & r1945 & r1952 & r1953 & r1954 & r1955 & r1962 & r1963 & r1964 & r1965);
        r1793 := r1973;
      end if;
      r1660 := r1793;
    end if;
    return r1660;
  end rewire_expwords_1657;
  function rewire_littleendianp_1695(r1696 : std_logic_vector) return std_logic_vector
  is
    variable r1774 : std_logic_vector(0 to 31) := (others => '0');
    variable r1773 : std_logic_vector(0 to 7) := (others => '0');
    variable r1771 : std_logic_vector(0 to 7) := (others => '0');
    variable r1769 : std_logic_vector(0 to 7) := (others => '0');
    variable r1767 : std_logic_vector(0 to 7) := (others => '0');
    variable EMPTY : std_logic_vector(0 to -1) := (others => '0');
    variable b1764 : boolean := false;
    variable b1763 : boolean := false;
    variable b1762 : boolean := false;
    variable b1761 : boolean := false;
    variable b1760 : boolean := false;
    variable b1759 : boolean := false;
    variable b1758 : boolean := false;
    variable b1757 : boolean := false;
    variable b1756 : boolean := false;
    variable b1755 : boolean := false;
    variable b1754 : boolean := false;
    variable b1753 : boolean := false;
    variable b1752 : boolean := false;
    variable b1751 : boolean := false;
    variable b1750 : boolean := false;
    variable b1749 : boolean := false;
    variable b1748 : boolean := false;
    variable b1747 : boolean := false;
    variable b1746 : boolean := false;
    variable b1745 : boolean := false;
    variable b1744 : boolean := false;
    variable b1743 : boolean := false;
    variable b1742 : boolean := false;
    variable b1741 : boolean := false;
    variable b1740 : boolean := false;
    variable b1739 : boolean := false;
    variable b1738 : boolean := false;
    variable b1737 : boolean := false;
    variable b1736 : boolean := false;
    variable b1735 : boolean := false;
    variable b1734 : boolean := false;
    variable b1733 : boolean := false;
    variable b1732 : boolean := false;
    variable r1731 : std_logic_vector(0 to 0) := (others => '0');
    variable r1730 : std_logic_vector(0 to 0) := (others => '0');
    variable r1729 : std_logic_vector(0 to 0) := (others => '0');
    variable r1728 : std_logic_vector(0 to 0) := (others => '0');
    variable r1727 : std_logic_vector(0 to 0) := (others => '0');
    variable r1726 : std_logic_vector(0 to 0) := (others => '0');
    variable r1725 : std_logic_vector(0 to 0) := (others => '0');
    variable r1724 : std_logic_vector(0 to 0) := (others => '0');
    variable r1723 : std_logic_vector(0 to 0) := (others => '0');
    variable r1722 : std_logic_vector(0 to 0) := (others => '0');
    variable r1721 : std_logic_vector(0 to 0) := (others => '0');
    variable r1720 : std_logic_vector(0 to 0) := (others => '0');
    variable r1719 : std_logic_vector(0 to 0) := (others => '0');
    variable r1718 : std_logic_vector(0 to 0) := (others => '0');
    variable r1717 : std_logic_vector(0 to 0) := (others => '0');
    variable r1716 : std_logic_vector(0 to 0) := (others => '0');
    variable r1715 : std_logic_vector(0 to 0) := (others => '0');
    variable r1714 : std_logic_vector(0 to 0) := (others => '0');
    variable r1713 : std_logic_vector(0 to 0) := (others => '0');
    variable r1712 : std_logic_vector(0 to 0) := (others => '0');
    variable r1711 : std_logic_vector(0 to 0) := (others => '0');
    variable r1710 : std_logic_vector(0 to 0) := (others => '0');
    variable r1709 : std_logic_vector(0 to 0) := (others => '0');
    variable r1708 : std_logic_vector(0 to 0) := (others => '0');
    variable r1707 : std_logic_vector(0 to 0) := (others => '0');
    variable r1706 : std_logic_vector(0 to 0) := (others => '0');
    variable r1705 : std_logic_vector(0 to 0) := (others => '0');
    variable r1704 : std_logic_vector(0 to 0) := (others => '0');
    variable r1703 : std_logic_vector(0 to 0) := (others => '0');
    variable r1702 : std_logic_vector(0 to 0) := (others => '0');
    variable r1701 : std_logic_vector(0 to 0) := (others => '0');
    variable r1700 : std_logic_vector(0 to 0) := (others => '0');
    variable b1699 : boolean := false;
    variable r1698 : std_logic_vector(0 to 31) := (others => '0');
  begin
    b1699 := true;
    r1700 := r1696(0 to 0);
    r1701 := r1696(1 to 1);
    r1702 := r1696(2 to 2);
    r1703 := r1696(3 to 3);
    r1704 := r1696(4 to 4);
    r1705 := r1696(5 to 5);
    r1706 := r1696(6 to 6);
    r1707 := r1696(7 to 7);
    r1708 := r1696(8 to 8);
    r1709 := r1696(9 to 9);
    r1710 := r1696(10 to 10);
    r1711 := r1696(11 to 11);
    r1712 := r1696(12 to 12);
    r1713 := r1696(13 to 13);
    r1714 := r1696(14 to 14);
    r1715 := r1696(15 to 15);
    r1716 := r1696(16 to 16);
    r1717 := r1696(17 to 17);
    r1718 := r1696(18 to 18);
    r1719 := r1696(19 to 19);
    r1720 := r1696(20 to 20);
    r1721 := r1696(21 to 21);
    r1722 := r1696(22 to 22);
    r1723 := r1696(23 to 23);
    r1724 := r1696(24 to 24);
    r1725 := r1696(25 to 25);
    r1726 := r1696(26 to 26);
    r1727 := r1696(27 to 27);
    r1728 := r1696(28 to 28);
    r1729 := r1696(29 to 29);
    r1730 := r1696(30 to 30);
    r1731 := r1696(31 to 31);
    b1732 := true;
    b1733 := true;
    b1734 := true;
    b1735 := true;
    b1736 := true;
    b1737 := true;
    b1738 := true;
    b1739 := true;
    b1740 := true;
    b1741 := true;
    b1742 := true;
    b1743 := true;
    b1744 := true;
    b1745 := true;
    b1746 := true;
    b1747 := true;
    b1748 := true;
    b1749 := true;
    b1750 := true;
    b1751 := true;
    b1752 := true;
    b1753 := true;
    b1754 := true;
    b1755 := true;
    b1756 := true;
    b1757 := true;
    b1758 := true;
    b1759 := true;
    b1760 := true;
    b1761 := true;
    b1762 := true;
    b1763 := true;
    b1764 := (b1732 AND (b1733 AND (b1734 AND (b1735 AND (b1736 AND (b1737 AND (b1738 AND (b1739 AND (b1740 AND (b1741 AND (b1742 AND (b1743 AND (b1744 AND (b1745 AND (b1746 AND (b1747 AND (b1748 AND (b1749 AND (b1750 AND (b1751 AND (b1752 AND (b1753 AND (b1754 AND (b1755 AND (b1756 AND (b1757 AND (b1758 AND (b1759 AND (b1760 AND (b1761 AND (b1762 AND b1763)))))))))))))))))))))))))))))));
    if b1764 then
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      r1767 := (r1700 & r1701 & r1702 & r1703 & r1704 & r1705 & r1706 & r1707);
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      r1769 := (r1708 & r1709 & r1710 & r1711 & r1712 & r1713 & r1714 & r1715);
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      r1771 := (r1716 & r1717 & r1718 & r1719 & r1720 & r1721 & r1722 & r1723);
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      r1773 := (r1724 & r1725 & r1726 & r1727 & r1728 & r1729 & r1730 & r1731);
      r1774 := (r1767 & r1769 & r1771 & r1773);
      r1698 := r1774;
    end if;
    return r1698;
  end rewire_littleendianp_1695;
  function rewire_sigma3_1529 return std_logic_vector
  is
    variable r1604 : std_logic_vector(0 to 31) := (others => '0');
    variable r1603 : std_logic_vector(0 to 7) := (others => '0');
    variable r1601 : std_logic_vector(0 to 0) := (others => '0');
    variable r1599 : std_logic_vector(0 to 0) := (others => '0');
    variable r1597 : std_logic_vector(0 to 0) := (others => '0');
    variable r1595 : std_logic_vector(0 to 0) := (others => '0');
    variable r1593 : std_logic_vector(0 to 0) := (others => '0');
    variable r1591 : std_logic_vector(0 to 0) := (others => '0');
    variable r1589 : std_logic_vector(0 to 0) := (others => '0');
    variable r1587 : std_logic_vector(0 to 0) := (others => '0');
    variable r1585 : std_logic_vector(0 to 7) := (others => '0');
    variable r1583 : std_logic_vector(0 to 0) := (others => '0');
    variable r1581 : std_logic_vector(0 to 0) := (others => '0');
    variable r1579 : std_logic_vector(0 to 0) := (others => '0');
    variable r1577 : std_logic_vector(0 to 0) := (others => '0');
    variable r1575 : std_logic_vector(0 to 0) := (others => '0');
    variable r1573 : std_logic_vector(0 to 0) := (others => '0');
    variable r1571 : std_logic_vector(0 to 0) := (others => '0');
    variable r1569 : std_logic_vector(0 to 0) := (others => '0');
    variable r1567 : std_logic_vector(0 to 7) := (others => '0');
    variable r1565 : std_logic_vector(0 to 0) := (others => '0');
    variable r1563 : std_logic_vector(0 to 0) := (others => '0');
    variable r1561 : std_logic_vector(0 to 0) := (others => '0');
    variable r1559 : std_logic_vector(0 to 0) := (others => '0');
    variable r1557 : std_logic_vector(0 to 0) := (others => '0');
    variable r1555 : std_logic_vector(0 to 0) := (others => '0');
    variable r1553 : std_logic_vector(0 to 0) := (others => '0');
    variable r1551 : std_logic_vector(0 to 0) := (others => '0');
    variable r1549 : std_logic_vector(0 to 7) := (others => '0');
    variable r1547 : std_logic_vector(0 to 0) := (others => '0');
    variable r1545 : std_logic_vector(0 to 0) := (others => '0');
    variable r1543 : std_logic_vector(0 to 0) := (others => '0');
    variable r1541 : std_logic_vector(0 to 0) := (others => '0');
    variable r1539 : std_logic_vector(0 to 0) := (others => '0');
    variable r1537 : std_logic_vector(0 to 0) := (others => '0');
    variable r1535 : std_logic_vector(0 to 0) := (others => '0');
    variable r1533 : std_logic_vector(0 to 0) := (others => '0');
    variable EMPTY : std_logic_vector(0 to -1) := (others => '0');
  begin
    r1533 := "0";
    r1535 := "0";
    r1537 := "1";
    r1539 := "0";
    r1541 := "1";
    r1543 := "1";
    r1545 := "1";
    r1547 := "0";
    r1549 := (r1533 & r1535 & r1537 & r1539 & r1541 & r1543 & r1545 & r1547);
    r1551 := "1";
    r1553 := "0";
    r1555 := "1";
    r1557 := "0";
    r1559 := "0";
    r1561 := "1";
    r1563 := "1";
    r1565 := "0";
    r1567 := (r1551 & r1553 & r1555 & r1557 & r1559 & r1561 & r1563 & r1565);
    r1569 := "0";
    r1571 := "0";
    r1573 := "0";
    r1575 := "0";
    r1577 := "0";
    r1579 := "1";
    r1581 := "0";
    r1583 := "0";
    r1585 := (r1569 & r1571 & r1573 & r1575 & r1577 & r1579 & r1581 & r1583);
    r1587 := "1";
    r1589 := "1";
    r1591 := "0";
    r1593 := "1";
    r1595 := "0";
    r1597 := "1";
    r1599 := "1";
    r1601 := "0";
    r1603 := (r1587 & r1589 & r1591 & r1593 & r1595 & r1597 & r1599 & r1601);
    r1604 := (r1549 & r1567 & r1585 & r1603);
    return r1604;
  end rewire_sigma3_1529;
  function rewire_sigma2_1452 return std_logic_vector
  is
    variable r1527 : std_logic_vector(0 to 31) := (others => '0');
    variable r1526 : std_logic_vector(0 to 7) := (others => '0');
    variable r1524 : std_logic_vector(0 to 0) := (others => '0');
    variable r1522 : std_logic_vector(0 to 0) := (others => '0');
    variable r1520 : std_logic_vector(0 to 0) := (others => '0');
    variable r1518 : std_logic_vector(0 to 0) := (others => '0');
    variable r1516 : std_logic_vector(0 to 0) := (others => '0');
    variable r1514 : std_logic_vector(0 to 0) := (others => '0');
    variable r1512 : std_logic_vector(0 to 0) := (others => '0');
    variable r1510 : std_logic_vector(0 to 0) := (others => '0');
    variable r1508 : std_logic_vector(0 to 7) := (others => '0');
    variable r1506 : std_logic_vector(0 to 0) := (others => '0');
    variable r1504 : std_logic_vector(0 to 0) := (others => '0');
    variable r1502 : std_logic_vector(0 to 0) := (others => '0');
    variable r1500 : std_logic_vector(0 to 0) := (others => '0');
    variable r1498 : std_logic_vector(0 to 0) := (others => '0');
    variable r1496 : std_logic_vector(0 to 0) := (others => '0');
    variable r1494 : std_logic_vector(0 to 0) := (others => '0');
    variable r1492 : std_logic_vector(0 to 0) := (others => '0');
    variable r1490 : std_logic_vector(0 to 7) := (others => '0');
    variable r1488 : std_logic_vector(0 to 0) := (others => '0');
    variable r1486 : std_logic_vector(0 to 0) := (others => '0');
    variable r1484 : std_logic_vector(0 to 0) := (others => '0');
    variable r1482 : std_logic_vector(0 to 0) := (others => '0');
    variable r1480 : std_logic_vector(0 to 0) := (others => '0');
    variable r1478 : std_logic_vector(0 to 0) := (others => '0');
    variable r1476 : std_logic_vector(0 to 0) := (others => '0');
    variable r1474 : std_logic_vector(0 to 0) := (others => '0');
    variable r1472 : std_logic_vector(0 to 7) := (others => '0');
    variable r1470 : std_logic_vector(0 to 0) := (others => '0');
    variable r1468 : std_logic_vector(0 to 0) := (others => '0');
    variable r1466 : std_logic_vector(0 to 0) := (others => '0');
    variable r1464 : std_logic_vector(0 to 0) := (others => '0');
    variable r1462 : std_logic_vector(0 to 0) := (others => '0');
    variable r1460 : std_logic_vector(0 to 0) := (others => '0');
    variable r1458 : std_logic_vector(0 to 0) := (others => '0');
    variable r1456 : std_logic_vector(0 to 0) := (others => '0');
    variable EMPTY : std_logic_vector(0 to -1) := (others => '0');
  begin
    r1456 := "0";
    r1458 := "1";
    r1460 := "0";
    r1462 := "0";
    r1464 := "1";
    r1466 := "1";
    r1468 := "0";
    r1470 := "0";
    r1472 := (r1456 & r1458 & r1460 & r1462 & r1464 & r1466 & r1468 & r1470);
    r1474 := "1";
    r1476 := "0";
    r1478 := "1";
    r1480 := "1";
    r1482 := "0";
    r1484 := "1";
    r1486 := "0";
    r1488 := "0";
    r1490 := (r1474 & r1476 & r1478 & r1480 & r1482 & r1484 & r1486 & r1488);
    r1492 := "0";
    r1494 := "1";
    r1496 := "0";
    r1498 := "0";
    r1500 := "0";
    r1502 := "1";
    r1504 := "1";
    r1506 := "0";
    r1508 := (r1492 & r1494 & r1496 & r1498 & r1500 & r1502 & r1504 & r1506);
    r1510 := "1";
    r1512 := "0";
    r1514 := "0";
    r1516 := "1";
    r1518 := "1";
    r1520 := "1";
    r1522 := "1";
    r1524 := "0";
    r1526 := (r1510 & r1512 & r1514 & r1516 & r1518 & r1520 & r1522 & r1524);
    r1527 := (r1472 & r1490 & r1508 & r1526);
    return r1527;
  end rewire_sigma2_1452;
  function rewire_sigma1_1375 return std_logic_vector
  is
    variable r1450 : std_logic_vector(0 to 31) := (others => '0');
    variable r1449 : std_logic_vector(0 to 7) := (others => '0');
    variable r1447 : std_logic_vector(0 to 0) := (others => '0');
    variable r1445 : std_logic_vector(0 to 0) := (others => '0');
    variable r1443 : std_logic_vector(0 to 0) := (others => '0');
    variable r1441 : std_logic_vector(0 to 0) := (others => '0');
    variable r1439 : std_logic_vector(0 to 0) := (others => '0');
    variable r1437 : std_logic_vector(0 to 0) := (others => '0');
    variable r1435 : std_logic_vector(0 to 0) := (others => '0');
    variable r1433 : std_logic_vector(0 to 0) := (others => '0');
    variable r1431 : std_logic_vector(0 to 7) := (others => '0');
    variable r1429 : std_logic_vector(0 to 0) := (others => '0');
    variable r1427 : std_logic_vector(0 to 0) := (others => '0');
    variable r1425 : std_logic_vector(0 to 0) := (others => '0');
    variable r1423 : std_logic_vector(0 to 0) := (others => '0');
    variable r1421 : std_logic_vector(0 to 0) := (others => '0');
    variable r1419 : std_logic_vector(0 to 0) := (others => '0');
    variable r1417 : std_logic_vector(0 to 0) := (others => '0');
    variable r1415 : std_logic_vector(0 to 0) := (others => '0');
    variable r1413 : std_logic_vector(0 to 7) := (others => '0');
    variable r1411 : std_logic_vector(0 to 0) := (others => '0');
    variable r1409 : std_logic_vector(0 to 0) := (others => '0');
    variable r1407 : std_logic_vector(0 to 0) := (others => '0');
    variable r1405 : std_logic_vector(0 to 0) := (others => '0');
    variable r1403 : std_logic_vector(0 to 0) := (others => '0');
    variable r1401 : std_logic_vector(0 to 0) := (others => '0');
    variable r1399 : std_logic_vector(0 to 0) := (others => '0');
    variable r1397 : std_logic_vector(0 to 0) := (others => '0');
    variable r1395 : std_logic_vector(0 to 7) := (others => '0');
    variable r1393 : std_logic_vector(0 to 0) := (others => '0');
    variable r1391 : std_logic_vector(0 to 0) := (others => '0');
    variable r1389 : std_logic_vector(0 to 0) := (others => '0');
    variable r1387 : std_logic_vector(0 to 0) := (others => '0');
    variable r1385 : std_logic_vector(0 to 0) := (others => '0');
    variable r1383 : std_logic_vector(0 to 0) := (others => '0');
    variable r1381 : std_logic_vector(0 to 0) := (others => '0');
    variable r1379 : std_logic_vector(0 to 0) := (others => '0');
    variable EMPTY : std_logic_vector(0 to -1) := (others => '0');
  begin
    r1379 := "0";
    r1381 := "1";
    r1383 := "1";
    r1385 := "1";
    r1387 := "0";
    r1389 := "1";
    r1391 := "1";
    r1393 := "0";
    r1395 := (r1379 & r1381 & r1383 & r1385 & r1387 & r1389 & r1391 & r1393);
    r1397 := "0";
    r1399 := "0";
    r1401 := "1";
    r1403 := "0";
    r1405 := "0";
    r1407 := "1";
    r1409 := "1";
    r1411 := "0";
    r1413 := (r1397 & r1399 & r1401 & r1403 & r1405 & r1407 & r1409 & r1411);
    r1415 := "0";
    r1417 := "0";
    r1419 := "0";
    r1421 := "0";
    r1423 := "0";
    r1425 := "1";
    r1427 := "0";
    r1429 := "0";
    r1431 := (r1415 & r1417 & r1419 & r1421 & r1423 & r1425 & r1427 & r1429);
    r1433 := "1";
    r1435 := "1";
    r1437 := "0";
    r1439 := "0";
    r1441 := "1";
    r1443 := "1";
    r1445 := "0";
    r1447 := "0";
    r1449 := (r1433 & r1435 & r1437 & r1439 & r1441 & r1443 & r1445 & r1447);
    r1450 := (r1395 & r1413 & r1431 & r1449);
    return r1450;
  end rewire_sigma1_1375;
  function rewire_sigma0_1298 return std_logic_vector
  is
    variable r1373 : std_logic_vector(0 to 31) := (others => '0');
    variable r1372 : std_logic_vector(0 to 7) := (others => '0');
    variable r1370 : std_logic_vector(0 to 0) := (others => '0');
    variable r1368 : std_logic_vector(0 to 0) := (others => '0');
    variable r1366 : std_logic_vector(0 to 0) := (others => '0');
    variable r1364 : std_logic_vector(0 to 0) := (others => '0');
    variable r1362 : std_logic_vector(0 to 0) := (others => '0');
    variable r1360 : std_logic_vector(0 to 0) := (others => '0');
    variable r1358 : std_logic_vector(0 to 0) := (others => '0');
    variable r1356 : std_logic_vector(0 to 0) := (others => '0');
    variable r1354 : std_logic_vector(0 to 7) := (others => '0');
    variable r1352 : std_logic_vector(0 to 0) := (others => '0');
    variable r1350 : std_logic_vector(0 to 0) := (others => '0');
    variable r1348 : std_logic_vector(0 to 0) := (others => '0');
    variable r1346 : std_logic_vector(0 to 0) := (others => '0');
    variable r1344 : std_logic_vector(0 to 0) := (others => '0');
    variable r1342 : std_logic_vector(0 to 0) := (others => '0');
    variable r1340 : std_logic_vector(0 to 0) := (others => '0');
    variable r1338 : std_logic_vector(0 to 0) := (others => '0');
    variable r1336 : std_logic_vector(0 to 7) := (others => '0');
    variable r1334 : std_logic_vector(0 to 0) := (others => '0');
    variable r1332 : std_logic_vector(0 to 0) := (others => '0');
    variable r1330 : std_logic_vector(0 to 0) := (others => '0');
    variable r1328 : std_logic_vector(0 to 0) := (others => '0');
    variable r1326 : std_logic_vector(0 to 0) := (others => '0');
    variable r1324 : std_logic_vector(0 to 0) := (others => '0');
    variable r1322 : std_logic_vector(0 to 0) := (others => '0');
    variable r1320 : std_logic_vector(0 to 0) := (others => '0');
    variable r1318 : std_logic_vector(0 to 7) := (others => '0');
    variable r1316 : std_logic_vector(0 to 0) := (others => '0');
    variable r1314 : std_logic_vector(0 to 0) := (others => '0');
    variable r1312 : std_logic_vector(0 to 0) := (others => '0');
    variable r1310 : std_logic_vector(0 to 0) := (others => '0');
    variable r1308 : std_logic_vector(0 to 0) := (others => '0');
    variable r1306 : std_logic_vector(0 to 0) := (others => '0');
    variable r1304 : std_logic_vector(0 to 0) := (others => '0');
    variable r1302 : std_logic_vector(0 to 0) := (others => '0');
    variable EMPTY : std_logic_vector(0 to -1) := (others => '0');
  begin
    r1302 := "1";
    r1304 := "0";
    r1306 := "1";
    r1308 := "0";
    r1310 := "0";
    r1312 := "1";
    r1314 := "1";
    r1316 := "0";
    r1318 := (r1302 & r1304 & r1306 & r1308 & r1310 & r1312 & r1314 & r1316);
    r1320 := "0";
    r1322 := "0";
    r1324 := "0";
    r1326 := "1";
    r1328 := "1";
    r1330 := "1";
    r1332 := "1";
    r1334 := "0";
    r1336 := (r1320 & r1322 & r1324 & r1326 & r1328 & r1330 & r1332 & r1334);
    r1338 := "0";
    r1340 := "0";
    r1342 := "0";
    r1344 := "0";
    r1346 := "1";
    r1348 := "1";
    r1350 := "1";
    r1352 := "0";
    r1354 := (r1338 & r1340 & r1342 & r1344 & r1346 & r1348 & r1350 & r1352);
    r1356 := "1";
    r1358 := "0";
    r1360 := "0";
    r1362 := "0";
    r1364 := "0";
    r1366 := "1";
    r1368 := "1";
    r1370 := "0";
    r1372 := (r1356 & r1358 & r1360 & r1362 & r1364 & r1366 & r1368 & r1370);
    r1373 := (r1318 & r1336 & r1354 & r1372);
    return r1373;
  end rewire_sigma0_1298;
  function rewire_zerothoutput_3 return std_logic_vector
  is
    variable r1158 : std_logic_vector(0 to 511) := (others => '0');
    variable r1157 : std_logic_vector(0 to 7) := (others => '0');
    variable r1155 : std_logic_vector(0 to 0) := (others => '0');
    variable r1153 : std_logic_vector(0 to 0) := (others => '0');
    variable r1151 : std_logic_vector(0 to 0) := (others => '0');
    variable r1149 : std_logic_vector(0 to 0) := (others => '0');
    variable r1147 : std_logic_vector(0 to 0) := (others => '0');
    variable r1145 : std_logic_vector(0 to 0) := (others => '0');
    variable r1143 : std_logic_vector(0 to 0) := (others => '0');
    variable r1141 : std_logic_vector(0 to 0) := (others => '0');
    variable r1139 : std_logic_vector(0 to 7) := (others => '0');
    variable r1137 : std_logic_vector(0 to 0) := (others => '0');
    variable r1135 : std_logic_vector(0 to 0) := (others => '0');
    variable r1133 : std_logic_vector(0 to 0) := (others => '0');
    variable r1131 : std_logic_vector(0 to 0) := (others => '0');
    variable r1129 : std_logic_vector(0 to 0) := (others => '0');
    variable r1127 : std_logic_vector(0 to 0) := (others => '0');
    variable r1125 : std_logic_vector(0 to 0) := (others => '0');
    variable r1123 : std_logic_vector(0 to 0) := (others => '0');
    variable r1121 : std_logic_vector(0 to 7) := (others => '0');
    variable r1119 : std_logic_vector(0 to 0) := (others => '0');
    variable r1117 : std_logic_vector(0 to 0) := (others => '0');
    variable r1115 : std_logic_vector(0 to 0) := (others => '0');
    variable r1113 : std_logic_vector(0 to 0) := (others => '0');
    variable r1111 : std_logic_vector(0 to 0) := (others => '0');
    variable r1109 : std_logic_vector(0 to 0) := (others => '0');
    variable r1107 : std_logic_vector(0 to 0) := (others => '0');
    variable r1105 : std_logic_vector(0 to 0) := (others => '0');
    variable r1103 : std_logic_vector(0 to 7) := (others => '0');
    variable r1101 : std_logic_vector(0 to 0) := (others => '0');
    variable r1099 : std_logic_vector(0 to 0) := (others => '0');
    variable r1097 : std_logic_vector(0 to 0) := (others => '0');
    variable r1095 : std_logic_vector(0 to 0) := (others => '0');
    variable r1093 : std_logic_vector(0 to 0) := (others => '0');
    variable r1091 : std_logic_vector(0 to 0) := (others => '0');
    variable r1089 : std_logic_vector(0 to 0) := (others => '0');
    variable r1087 : std_logic_vector(0 to 0) := (others => '0');
    variable r1085 : std_logic_vector(0 to 7) := (others => '0');
    variable r1083 : std_logic_vector(0 to 0) := (others => '0');
    variable r1081 : std_logic_vector(0 to 0) := (others => '0');
    variable r1079 : std_logic_vector(0 to 0) := (others => '0');
    variable r1077 : std_logic_vector(0 to 0) := (others => '0');
    variable r1075 : std_logic_vector(0 to 0) := (others => '0');
    variable r1073 : std_logic_vector(0 to 0) := (others => '0');
    variable r1071 : std_logic_vector(0 to 0) := (others => '0');
    variable r1069 : std_logic_vector(0 to 0) := (others => '0');
    variable r1067 : std_logic_vector(0 to 7) := (others => '0');
    variable r1065 : std_logic_vector(0 to 0) := (others => '0');
    variable r1063 : std_logic_vector(0 to 0) := (others => '0');
    variable r1061 : std_logic_vector(0 to 0) := (others => '0');
    variable r1059 : std_logic_vector(0 to 0) := (others => '0');
    variable r1057 : std_logic_vector(0 to 0) := (others => '0');
    variable r1055 : std_logic_vector(0 to 0) := (others => '0');
    variable r1053 : std_logic_vector(0 to 0) := (others => '0');
    variable r1051 : std_logic_vector(0 to 0) := (others => '0');
    variable r1049 : std_logic_vector(0 to 7) := (others => '0');
    variable r1047 : std_logic_vector(0 to 0) := (others => '0');
    variable r1045 : std_logic_vector(0 to 0) := (others => '0');
    variable r1043 : std_logic_vector(0 to 0) := (others => '0');
    variable r1041 : std_logic_vector(0 to 0) := (others => '0');
    variable r1039 : std_logic_vector(0 to 0) := (others => '0');
    variable r1037 : std_logic_vector(0 to 0) := (others => '0');
    variable r1035 : std_logic_vector(0 to 0) := (others => '0');
    variable r1033 : std_logic_vector(0 to 0) := (others => '0');
    variable r1031 : std_logic_vector(0 to 7) := (others => '0');
    variable r1029 : std_logic_vector(0 to 0) := (others => '0');
    variable r1027 : std_logic_vector(0 to 0) := (others => '0');
    variable r1025 : std_logic_vector(0 to 0) := (others => '0');
    variable r1023 : std_logic_vector(0 to 0) := (others => '0');
    variable r1021 : std_logic_vector(0 to 0) := (others => '0');
    variable r1019 : std_logic_vector(0 to 0) := (others => '0');
    variable r1017 : std_logic_vector(0 to 0) := (others => '0');
    variable r1015 : std_logic_vector(0 to 0) := (others => '0');
    variable r1013 : std_logic_vector(0 to 7) := (others => '0');
    variable r1011 : std_logic_vector(0 to 0) := (others => '0');
    variable r1009 : std_logic_vector(0 to 0) := (others => '0');
    variable r1007 : std_logic_vector(0 to 0) := (others => '0');
    variable r1005 : std_logic_vector(0 to 0) := (others => '0');
    variable r1003 : std_logic_vector(0 to 0) := (others => '0');
    variable r1001 : std_logic_vector(0 to 0) := (others => '0');
    variable r999 : std_logic_vector(0 to 0) := (others => '0');
    variable r997 : std_logic_vector(0 to 0) := (others => '0');
    variable r995 : std_logic_vector(0 to 7) := (others => '0');
    variable r993 : std_logic_vector(0 to 0) := (others => '0');
    variable r991 : std_logic_vector(0 to 0) := (others => '0');
    variable r989 : std_logic_vector(0 to 0) := (others => '0');
    variable r987 : std_logic_vector(0 to 0) := (others => '0');
    variable r985 : std_logic_vector(0 to 0) := (others => '0');
    variable r983 : std_logic_vector(0 to 0) := (others => '0');
    variable r981 : std_logic_vector(0 to 0) := (others => '0');
    variable r979 : std_logic_vector(0 to 0) := (others => '0');
    variable r977 : std_logic_vector(0 to 7) := (others => '0');
    variable r975 : std_logic_vector(0 to 0) := (others => '0');
    variable r973 : std_logic_vector(0 to 0) := (others => '0');
    variable r971 : std_logic_vector(0 to 0) := (others => '0');
    variable r969 : std_logic_vector(0 to 0) := (others => '0');
    variable r967 : std_logic_vector(0 to 0) := (others => '0');
    variable r965 : std_logic_vector(0 to 0) := (others => '0');
    variable r963 : std_logic_vector(0 to 0) := (others => '0');
    variable r961 : std_logic_vector(0 to 0) := (others => '0');
    variable r959 : std_logic_vector(0 to 7) := (others => '0');
    variable r957 : std_logic_vector(0 to 0) := (others => '0');
    variable r955 : std_logic_vector(0 to 0) := (others => '0');
    variable r953 : std_logic_vector(0 to 0) := (others => '0');
    variable r951 : std_logic_vector(0 to 0) := (others => '0');
    variable r949 : std_logic_vector(0 to 0) := (others => '0');
    variable r947 : std_logic_vector(0 to 0) := (others => '0');
    variable r945 : std_logic_vector(0 to 0) := (others => '0');
    variable r943 : std_logic_vector(0 to 0) := (others => '0');
    variable r941 : std_logic_vector(0 to 7) := (others => '0');
    variable r939 : std_logic_vector(0 to 0) := (others => '0');
    variable r937 : std_logic_vector(0 to 0) := (others => '0');
    variable r935 : std_logic_vector(0 to 0) := (others => '0');
    variable r933 : std_logic_vector(0 to 0) := (others => '0');
    variable r931 : std_logic_vector(0 to 0) := (others => '0');
    variable r929 : std_logic_vector(0 to 0) := (others => '0');
    variable r927 : std_logic_vector(0 to 0) := (others => '0');
    variable r925 : std_logic_vector(0 to 0) := (others => '0');
    variable r923 : std_logic_vector(0 to 7) := (others => '0');
    variable r921 : std_logic_vector(0 to 0) := (others => '0');
    variable r919 : std_logic_vector(0 to 0) := (others => '0');
    variable r917 : std_logic_vector(0 to 0) := (others => '0');
    variable r915 : std_logic_vector(0 to 0) := (others => '0');
    variable r913 : std_logic_vector(0 to 0) := (others => '0');
    variable r911 : std_logic_vector(0 to 0) := (others => '0');
    variable r909 : std_logic_vector(0 to 0) := (others => '0');
    variable r907 : std_logic_vector(0 to 0) := (others => '0');
    variable r905 : std_logic_vector(0 to 7) := (others => '0');
    variable r903 : std_logic_vector(0 to 0) := (others => '0');
    variable r901 : std_logic_vector(0 to 0) := (others => '0');
    variable r899 : std_logic_vector(0 to 0) := (others => '0');
    variable r897 : std_logic_vector(0 to 0) := (others => '0');
    variable r895 : std_logic_vector(0 to 0) := (others => '0');
    variable r893 : std_logic_vector(0 to 0) := (others => '0');
    variable r891 : std_logic_vector(0 to 0) := (others => '0');
    variable r889 : std_logic_vector(0 to 0) := (others => '0');
    variable r887 : std_logic_vector(0 to 7) := (others => '0');
    variable r885 : std_logic_vector(0 to 0) := (others => '0');
    variable r883 : std_logic_vector(0 to 0) := (others => '0');
    variable r881 : std_logic_vector(0 to 0) := (others => '0');
    variable r879 : std_logic_vector(0 to 0) := (others => '0');
    variable r877 : std_logic_vector(0 to 0) := (others => '0');
    variable r875 : std_logic_vector(0 to 0) := (others => '0');
    variable r873 : std_logic_vector(0 to 0) := (others => '0');
    variable r871 : std_logic_vector(0 to 0) := (others => '0');
    variable r869 : std_logic_vector(0 to 7) := (others => '0');
    variable r867 : std_logic_vector(0 to 0) := (others => '0');
    variable r865 : std_logic_vector(0 to 0) := (others => '0');
    variable r863 : std_logic_vector(0 to 0) := (others => '0');
    variable r861 : std_logic_vector(0 to 0) := (others => '0');
    variable r859 : std_logic_vector(0 to 0) := (others => '0');
    variable r857 : std_logic_vector(0 to 0) := (others => '0');
    variable r855 : std_logic_vector(0 to 0) := (others => '0');
    variable r853 : std_logic_vector(0 to 0) := (others => '0');
    variable r851 : std_logic_vector(0 to 7) := (others => '0');
    variable r849 : std_logic_vector(0 to 0) := (others => '0');
    variable r847 : std_logic_vector(0 to 0) := (others => '0');
    variable r845 : std_logic_vector(0 to 0) := (others => '0');
    variable r843 : std_logic_vector(0 to 0) := (others => '0');
    variable r841 : std_logic_vector(0 to 0) := (others => '0');
    variable r839 : std_logic_vector(0 to 0) := (others => '0');
    variable r837 : std_logic_vector(0 to 0) := (others => '0');
    variable r835 : std_logic_vector(0 to 0) := (others => '0');
    variable r833 : std_logic_vector(0 to 7) := (others => '0');
    variable r831 : std_logic_vector(0 to 0) := (others => '0');
    variable r829 : std_logic_vector(0 to 0) := (others => '0');
    variable r827 : std_logic_vector(0 to 0) := (others => '0');
    variable r825 : std_logic_vector(0 to 0) := (others => '0');
    variable r823 : std_logic_vector(0 to 0) := (others => '0');
    variable r821 : std_logic_vector(0 to 0) := (others => '0');
    variable r819 : std_logic_vector(0 to 0) := (others => '0');
    variable r817 : std_logic_vector(0 to 0) := (others => '0');
    variable r815 : std_logic_vector(0 to 7) := (others => '0');
    variable r813 : std_logic_vector(0 to 0) := (others => '0');
    variable r811 : std_logic_vector(0 to 0) := (others => '0');
    variable r809 : std_logic_vector(0 to 0) := (others => '0');
    variable r807 : std_logic_vector(0 to 0) := (others => '0');
    variable r805 : std_logic_vector(0 to 0) := (others => '0');
    variable r803 : std_logic_vector(0 to 0) := (others => '0');
    variable r801 : std_logic_vector(0 to 0) := (others => '0');
    variable r799 : std_logic_vector(0 to 0) := (others => '0');
    variable r797 : std_logic_vector(0 to 7) := (others => '0');
    variable r795 : std_logic_vector(0 to 0) := (others => '0');
    variable r793 : std_logic_vector(0 to 0) := (others => '0');
    variable r791 : std_logic_vector(0 to 0) := (others => '0');
    variable r789 : std_logic_vector(0 to 0) := (others => '0');
    variable r787 : std_logic_vector(0 to 0) := (others => '0');
    variable r785 : std_logic_vector(0 to 0) := (others => '0');
    variable r783 : std_logic_vector(0 to 0) := (others => '0');
    variable r781 : std_logic_vector(0 to 0) := (others => '0');
    variable r779 : std_logic_vector(0 to 7) := (others => '0');
    variable r777 : std_logic_vector(0 to 0) := (others => '0');
    variable r775 : std_logic_vector(0 to 0) := (others => '0');
    variable r773 : std_logic_vector(0 to 0) := (others => '0');
    variable r771 : std_logic_vector(0 to 0) := (others => '0');
    variable r769 : std_logic_vector(0 to 0) := (others => '0');
    variable r767 : std_logic_vector(0 to 0) := (others => '0');
    variable r765 : std_logic_vector(0 to 0) := (others => '0');
    variable r763 : std_logic_vector(0 to 0) := (others => '0');
    variable r761 : std_logic_vector(0 to 7) := (others => '0');
    variable r759 : std_logic_vector(0 to 0) := (others => '0');
    variable r757 : std_logic_vector(0 to 0) := (others => '0');
    variable r755 : std_logic_vector(0 to 0) := (others => '0');
    variable r753 : std_logic_vector(0 to 0) := (others => '0');
    variable r751 : std_logic_vector(0 to 0) := (others => '0');
    variable r749 : std_logic_vector(0 to 0) := (others => '0');
    variable r747 : std_logic_vector(0 to 0) := (others => '0');
    variable r745 : std_logic_vector(0 to 0) := (others => '0');
    variable r743 : std_logic_vector(0 to 7) := (others => '0');
    variable r741 : std_logic_vector(0 to 0) := (others => '0');
    variable r739 : std_logic_vector(0 to 0) := (others => '0');
    variable r737 : std_logic_vector(0 to 0) := (others => '0');
    variable r735 : std_logic_vector(0 to 0) := (others => '0');
    variable r733 : std_logic_vector(0 to 0) := (others => '0');
    variable r731 : std_logic_vector(0 to 0) := (others => '0');
    variable r729 : std_logic_vector(0 to 0) := (others => '0');
    variable r727 : std_logic_vector(0 to 0) := (others => '0');
    variable r725 : std_logic_vector(0 to 7) := (others => '0');
    variable r723 : std_logic_vector(0 to 0) := (others => '0');
    variable r721 : std_logic_vector(0 to 0) := (others => '0');
    variable r719 : std_logic_vector(0 to 0) := (others => '0');
    variable r717 : std_logic_vector(0 to 0) := (others => '0');
    variable r715 : std_logic_vector(0 to 0) := (others => '0');
    variable r713 : std_logic_vector(0 to 0) := (others => '0');
    variable r711 : std_logic_vector(0 to 0) := (others => '0');
    variable r709 : std_logic_vector(0 to 0) := (others => '0');
    variable r707 : std_logic_vector(0 to 7) := (others => '0');
    variable r705 : std_logic_vector(0 to 0) := (others => '0');
    variable r703 : std_logic_vector(0 to 0) := (others => '0');
    variable r701 : std_logic_vector(0 to 0) := (others => '0');
    variable r699 : std_logic_vector(0 to 0) := (others => '0');
    variable r697 : std_logic_vector(0 to 0) := (others => '0');
    variable r695 : std_logic_vector(0 to 0) := (others => '0');
    variable r693 : std_logic_vector(0 to 0) := (others => '0');
    variable r691 : std_logic_vector(0 to 0) := (others => '0');
    variable r689 : std_logic_vector(0 to 7) := (others => '0');
    variable r687 : std_logic_vector(0 to 0) := (others => '0');
    variable r685 : std_logic_vector(0 to 0) := (others => '0');
    variable r683 : std_logic_vector(0 to 0) := (others => '0');
    variable r681 : std_logic_vector(0 to 0) := (others => '0');
    variable r679 : std_logic_vector(0 to 0) := (others => '0');
    variable r677 : std_logic_vector(0 to 0) := (others => '0');
    variable r675 : std_logic_vector(0 to 0) := (others => '0');
    variable r673 : std_logic_vector(0 to 0) := (others => '0');
    variable r671 : std_logic_vector(0 to 7) := (others => '0');
    variable r669 : std_logic_vector(0 to 0) := (others => '0');
    variable r667 : std_logic_vector(0 to 0) := (others => '0');
    variable r665 : std_logic_vector(0 to 0) := (others => '0');
    variable r663 : std_logic_vector(0 to 0) := (others => '0');
    variable r661 : std_logic_vector(0 to 0) := (others => '0');
    variable r659 : std_logic_vector(0 to 0) := (others => '0');
    variable r657 : std_logic_vector(0 to 0) := (others => '0');
    variable r655 : std_logic_vector(0 to 0) := (others => '0');
    variable r653 : std_logic_vector(0 to 7) := (others => '0');
    variable r651 : std_logic_vector(0 to 0) := (others => '0');
    variable r649 : std_logic_vector(0 to 0) := (others => '0');
    variable r647 : std_logic_vector(0 to 0) := (others => '0');
    variable r645 : std_logic_vector(0 to 0) := (others => '0');
    variable r643 : std_logic_vector(0 to 0) := (others => '0');
    variable r641 : std_logic_vector(0 to 0) := (others => '0');
    variable r639 : std_logic_vector(0 to 0) := (others => '0');
    variable r637 : std_logic_vector(0 to 0) := (others => '0');
    variable r635 : std_logic_vector(0 to 7) := (others => '0');
    variable r633 : std_logic_vector(0 to 0) := (others => '0');
    variable r631 : std_logic_vector(0 to 0) := (others => '0');
    variable r629 : std_logic_vector(0 to 0) := (others => '0');
    variable r627 : std_logic_vector(0 to 0) := (others => '0');
    variable r625 : std_logic_vector(0 to 0) := (others => '0');
    variable r623 : std_logic_vector(0 to 0) := (others => '0');
    variable r621 : std_logic_vector(0 to 0) := (others => '0');
    variable r619 : std_logic_vector(0 to 0) := (others => '0');
    variable r617 : std_logic_vector(0 to 7) := (others => '0');
    variable r615 : std_logic_vector(0 to 0) := (others => '0');
    variable r613 : std_logic_vector(0 to 0) := (others => '0');
    variable r611 : std_logic_vector(0 to 0) := (others => '0');
    variable r609 : std_logic_vector(0 to 0) := (others => '0');
    variable r607 : std_logic_vector(0 to 0) := (others => '0');
    variable r605 : std_logic_vector(0 to 0) := (others => '0');
    variable r603 : std_logic_vector(0 to 0) := (others => '0');
    variable r601 : std_logic_vector(0 to 0) := (others => '0');
    variable r599 : std_logic_vector(0 to 7) := (others => '0');
    variable r597 : std_logic_vector(0 to 0) := (others => '0');
    variable r595 : std_logic_vector(0 to 0) := (others => '0');
    variable r593 : std_logic_vector(0 to 0) := (others => '0');
    variable r591 : std_logic_vector(0 to 0) := (others => '0');
    variable r589 : std_logic_vector(0 to 0) := (others => '0');
    variable r587 : std_logic_vector(0 to 0) := (others => '0');
    variable r585 : std_logic_vector(0 to 0) := (others => '0');
    variable r583 : std_logic_vector(0 to 0) := (others => '0');
    variable r581 : std_logic_vector(0 to 7) := (others => '0');
    variable r579 : std_logic_vector(0 to 0) := (others => '0');
    variable r577 : std_logic_vector(0 to 0) := (others => '0');
    variable r575 : std_logic_vector(0 to 0) := (others => '0');
    variable r573 : std_logic_vector(0 to 0) := (others => '0');
    variable r571 : std_logic_vector(0 to 0) := (others => '0');
    variable r569 : std_logic_vector(0 to 0) := (others => '0');
    variable r567 : std_logic_vector(0 to 0) := (others => '0');
    variable r565 : std_logic_vector(0 to 0) := (others => '0');
    variable r563 : std_logic_vector(0 to 7) := (others => '0');
    variable r561 : std_logic_vector(0 to 0) := (others => '0');
    variable r559 : std_logic_vector(0 to 0) := (others => '0');
    variable r557 : std_logic_vector(0 to 0) := (others => '0');
    variable r555 : std_logic_vector(0 to 0) := (others => '0');
    variable r553 : std_logic_vector(0 to 0) := (others => '0');
    variable r551 : std_logic_vector(0 to 0) := (others => '0');
    variable r549 : std_logic_vector(0 to 0) := (others => '0');
    variable r547 : std_logic_vector(0 to 0) := (others => '0');
    variable r545 : std_logic_vector(0 to 7) := (others => '0');
    variable r543 : std_logic_vector(0 to 0) := (others => '0');
    variable r541 : std_logic_vector(0 to 0) := (others => '0');
    variable r539 : std_logic_vector(0 to 0) := (others => '0');
    variable r537 : std_logic_vector(0 to 0) := (others => '0');
    variable r535 : std_logic_vector(0 to 0) := (others => '0');
    variable r533 : std_logic_vector(0 to 0) := (others => '0');
    variable r531 : std_logic_vector(0 to 0) := (others => '0');
    variable r529 : std_logic_vector(0 to 0) := (others => '0');
    variable r527 : std_logic_vector(0 to 7) := (others => '0');
    variable r525 : std_logic_vector(0 to 0) := (others => '0');
    variable r523 : std_logic_vector(0 to 0) := (others => '0');
    variable r521 : std_logic_vector(0 to 0) := (others => '0');
    variable r519 : std_logic_vector(0 to 0) := (others => '0');
    variable r517 : std_logic_vector(0 to 0) := (others => '0');
    variable r515 : std_logic_vector(0 to 0) := (others => '0');
    variable r513 : std_logic_vector(0 to 0) := (others => '0');
    variable r511 : std_logic_vector(0 to 0) := (others => '0');
    variable r509 : std_logic_vector(0 to 7) := (others => '0');
    variable r507 : std_logic_vector(0 to 0) := (others => '0');
    variable r505 : std_logic_vector(0 to 0) := (others => '0');
    variable r503 : std_logic_vector(0 to 0) := (others => '0');
    variable r501 : std_logic_vector(0 to 0) := (others => '0');
    variable r499 : std_logic_vector(0 to 0) := (others => '0');
    variable r497 : std_logic_vector(0 to 0) := (others => '0');
    variable r495 : std_logic_vector(0 to 0) := (others => '0');
    variable r493 : std_logic_vector(0 to 0) := (others => '0');
    variable r491 : std_logic_vector(0 to 7) := (others => '0');
    variable r489 : std_logic_vector(0 to 0) := (others => '0');
    variable r487 : std_logic_vector(0 to 0) := (others => '0');
    variable r485 : std_logic_vector(0 to 0) := (others => '0');
    variable r483 : std_logic_vector(0 to 0) := (others => '0');
    variable r481 : std_logic_vector(0 to 0) := (others => '0');
    variable r479 : std_logic_vector(0 to 0) := (others => '0');
    variable r477 : std_logic_vector(0 to 0) := (others => '0');
    variable r475 : std_logic_vector(0 to 0) := (others => '0');
    variable r473 : std_logic_vector(0 to 7) := (others => '0');
    variable r471 : std_logic_vector(0 to 0) := (others => '0');
    variable r469 : std_logic_vector(0 to 0) := (others => '0');
    variable r467 : std_logic_vector(0 to 0) := (others => '0');
    variable r465 : std_logic_vector(0 to 0) := (others => '0');
    variable r463 : std_logic_vector(0 to 0) := (others => '0');
    variable r461 : std_logic_vector(0 to 0) := (others => '0');
    variable r459 : std_logic_vector(0 to 0) := (others => '0');
    variable r457 : std_logic_vector(0 to 0) := (others => '0');
    variable r455 : std_logic_vector(0 to 7) := (others => '0');
    variable r453 : std_logic_vector(0 to 0) := (others => '0');
    variable r451 : std_logic_vector(0 to 0) := (others => '0');
    variable r449 : std_logic_vector(0 to 0) := (others => '0');
    variable r447 : std_logic_vector(0 to 0) := (others => '0');
    variable r445 : std_logic_vector(0 to 0) := (others => '0');
    variable r443 : std_logic_vector(0 to 0) := (others => '0');
    variable r441 : std_logic_vector(0 to 0) := (others => '0');
    variable r439 : std_logic_vector(0 to 0) := (others => '0');
    variable r437 : std_logic_vector(0 to 7) := (others => '0');
    variable r435 : std_logic_vector(0 to 0) := (others => '0');
    variable r433 : std_logic_vector(0 to 0) := (others => '0');
    variable r431 : std_logic_vector(0 to 0) := (others => '0');
    variable r429 : std_logic_vector(0 to 0) := (others => '0');
    variable r427 : std_logic_vector(0 to 0) := (others => '0');
    variable r425 : std_logic_vector(0 to 0) := (others => '0');
    variable r423 : std_logic_vector(0 to 0) := (others => '0');
    variable r421 : std_logic_vector(0 to 0) := (others => '0');
    variable r419 : std_logic_vector(0 to 7) := (others => '0');
    variable r417 : std_logic_vector(0 to 0) := (others => '0');
    variable r415 : std_logic_vector(0 to 0) := (others => '0');
    variable r413 : std_logic_vector(0 to 0) := (others => '0');
    variable r411 : std_logic_vector(0 to 0) := (others => '0');
    variable r409 : std_logic_vector(0 to 0) := (others => '0');
    variable r407 : std_logic_vector(0 to 0) := (others => '0');
    variable r405 : std_logic_vector(0 to 0) := (others => '0');
    variable r403 : std_logic_vector(0 to 0) := (others => '0');
    variable r401 : std_logic_vector(0 to 7) := (others => '0');
    variable r399 : std_logic_vector(0 to 0) := (others => '0');
    variable r397 : std_logic_vector(0 to 0) := (others => '0');
    variable r395 : std_logic_vector(0 to 0) := (others => '0');
    variable r393 : std_logic_vector(0 to 0) := (others => '0');
    variable r391 : std_logic_vector(0 to 0) := (others => '0');
    variable r389 : std_logic_vector(0 to 0) := (others => '0');
    variable r387 : std_logic_vector(0 to 0) := (others => '0');
    variable r385 : std_logic_vector(0 to 0) := (others => '0');
    variable r383 : std_logic_vector(0 to 7) := (others => '0');
    variable r381 : std_logic_vector(0 to 0) := (others => '0');
    variable r379 : std_logic_vector(0 to 0) := (others => '0');
    variable r377 : std_logic_vector(0 to 0) := (others => '0');
    variable r375 : std_logic_vector(0 to 0) := (others => '0');
    variable r373 : std_logic_vector(0 to 0) := (others => '0');
    variable r371 : std_logic_vector(0 to 0) := (others => '0');
    variable r369 : std_logic_vector(0 to 0) := (others => '0');
    variable r367 : std_logic_vector(0 to 0) := (others => '0');
    variable r365 : std_logic_vector(0 to 7) := (others => '0');
    variable r363 : std_logic_vector(0 to 0) := (others => '0');
    variable r361 : std_logic_vector(0 to 0) := (others => '0');
    variable r359 : std_logic_vector(0 to 0) := (others => '0');
    variable r357 : std_logic_vector(0 to 0) := (others => '0');
    variable r355 : std_logic_vector(0 to 0) := (others => '0');
    variable r353 : std_logic_vector(0 to 0) := (others => '0');
    variable r351 : std_logic_vector(0 to 0) := (others => '0');
    variable r349 : std_logic_vector(0 to 0) := (others => '0');
    variable r347 : std_logic_vector(0 to 7) := (others => '0');
    variable r345 : std_logic_vector(0 to 0) := (others => '0');
    variable r343 : std_logic_vector(0 to 0) := (others => '0');
    variable r341 : std_logic_vector(0 to 0) := (others => '0');
    variable r339 : std_logic_vector(0 to 0) := (others => '0');
    variable r337 : std_logic_vector(0 to 0) := (others => '0');
    variable r335 : std_logic_vector(0 to 0) := (others => '0');
    variable r333 : std_logic_vector(0 to 0) := (others => '0');
    variable r331 : std_logic_vector(0 to 0) := (others => '0');
    variable r329 : std_logic_vector(0 to 7) := (others => '0');
    variable r327 : std_logic_vector(0 to 0) := (others => '0');
    variable r325 : std_logic_vector(0 to 0) := (others => '0');
    variable r323 : std_logic_vector(0 to 0) := (others => '0');
    variable r321 : std_logic_vector(0 to 0) := (others => '0');
    variable r319 : std_logic_vector(0 to 0) := (others => '0');
    variable r317 : std_logic_vector(0 to 0) := (others => '0');
    variable r315 : std_logic_vector(0 to 0) := (others => '0');
    variable r313 : std_logic_vector(0 to 0) := (others => '0');
    variable r311 : std_logic_vector(0 to 7) := (others => '0');
    variable r309 : std_logic_vector(0 to 0) := (others => '0');
    variable r307 : std_logic_vector(0 to 0) := (others => '0');
    variable r305 : std_logic_vector(0 to 0) := (others => '0');
    variable r303 : std_logic_vector(0 to 0) := (others => '0');
    variable r301 : std_logic_vector(0 to 0) := (others => '0');
    variable r299 : std_logic_vector(0 to 0) := (others => '0');
    variable r297 : std_logic_vector(0 to 0) := (others => '0');
    variable r295 : std_logic_vector(0 to 0) := (others => '0');
    variable r293 : std_logic_vector(0 to 7) := (others => '0');
    variable r291 : std_logic_vector(0 to 0) := (others => '0');
    variable r289 : std_logic_vector(0 to 0) := (others => '0');
    variable r287 : std_logic_vector(0 to 0) := (others => '0');
    variable r285 : std_logic_vector(0 to 0) := (others => '0');
    variable r283 : std_logic_vector(0 to 0) := (others => '0');
    variable r281 : std_logic_vector(0 to 0) := (others => '0');
    variable r279 : std_logic_vector(0 to 0) := (others => '0');
    variable r277 : std_logic_vector(0 to 0) := (others => '0');
    variable r275 : std_logic_vector(0 to 7) := (others => '0');
    variable r273 : std_logic_vector(0 to 0) := (others => '0');
    variable r271 : std_logic_vector(0 to 0) := (others => '0');
    variable r269 : std_logic_vector(0 to 0) := (others => '0');
    variable r267 : std_logic_vector(0 to 0) := (others => '0');
    variable r265 : std_logic_vector(0 to 0) := (others => '0');
    variable r263 : std_logic_vector(0 to 0) := (others => '0');
    variable r261 : std_logic_vector(0 to 0) := (others => '0');
    variable r259 : std_logic_vector(0 to 0) := (others => '0');
    variable r257 : std_logic_vector(0 to 7) := (others => '0');
    variable r255 : std_logic_vector(0 to 0) := (others => '0');
    variable r253 : std_logic_vector(0 to 0) := (others => '0');
    variable r251 : std_logic_vector(0 to 0) := (others => '0');
    variable r249 : std_logic_vector(0 to 0) := (others => '0');
    variable r247 : std_logic_vector(0 to 0) := (others => '0');
    variable r245 : std_logic_vector(0 to 0) := (others => '0');
    variable r243 : std_logic_vector(0 to 0) := (others => '0');
    variable r241 : std_logic_vector(0 to 0) := (others => '0');
    variable r239 : std_logic_vector(0 to 7) := (others => '0');
    variable r237 : std_logic_vector(0 to 0) := (others => '0');
    variable r235 : std_logic_vector(0 to 0) := (others => '0');
    variable r233 : std_logic_vector(0 to 0) := (others => '0');
    variable r231 : std_logic_vector(0 to 0) := (others => '0');
    variable r229 : std_logic_vector(0 to 0) := (others => '0');
    variable r227 : std_logic_vector(0 to 0) := (others => '0');
    variable r225 : std_logic_vector(0 to 0) := (others => '0');
    variable r223 : std_logic_vector(0 to 0) := (others => '0');
    variable r221 : std_logic_vector(0 to 7) := (others => '0');
    variable r219 : std_logic_vector(0 to 0) := (others => '0');
    variable r217 : std_logic_vector(0 to 0) := (others => '0');
    variable r215 : std_logic_vector(0 to 0) := (others => '0');
    variable r213 : std_logic_vector(0 to 0) := (others => '0');
    variable r211 : std_logic_vector(0 to 0) := (others => '0');
    variable r209 : std_logic_vector(0 to 0) := (others => '0');
    variable r207 : std_logic_vector(0 to 0) := (others => '0');
    variable r205 : std_logic_vector(0 to 0) := (others => '0');
    variable r203 : std_logic_vector(0 to 7) := (others => '0');
    variable r201 : std_logic_vector(0 to 0) := (others => '0');
    variable r199 : std_logic_vector(0 to 0) := (others => '0');
    variable r197 : std_logic_vector(0 to 0) := (others => '0');
    variable r195 : std_logic_vector(0 to 0) := (others => '0');
    variable r193 : std_logic_vector(0 to 0) := (others => '0');
    variable r191 : std_logic_vector(0 to 0) := (others => '0');
    variable r189 : std_logic_vector(0 to 0) := (others => '0');
    variable r187 : std_logic_vector(0 to 0) := (others => '0');
    variable r185 : std_logic_vector(0 to 7) := (others => '0');
    variable r183 : std_logic_vector(0 to 0) := (others => '0');
    variable r181 : std_logic_vector(0 to 0) := (others => '0');
    variable r179 : std_logic_vector(0 to 0) := (others => '0');
    variable r177 : std_logic_vector(0 to 0) := (others => '0');
    variable r175 : std_logic_vector(0 to 0) := (others => '0');
    variable r173 : std_logic_vector(0 to 0) := (others => '0');
    variable r171 : std_logic_vector(0 to 0) := (others => '0');
    variable r169 : std_logic_vector(0 to 0) := (others => '0');
    variable r167 : std_logic_vector(0 to 7) := (others => '0');
    variable r165 : std_logic_vector(0 to 0) := (others => '0');
    variable r163 : std_logic_vector(0 to 0) := (others => '0');
    variable r161 : std_logic_vector(0 to 0) := (others => '0');
    variable r159 : std_logic_vector(0 to 0) := (others => '0');
    variable r157 : std_logic_vector(0 to 0) := (others => '0');
    variable r155 : std_logic_vector(0 to 0) := (others => '0');
    variable r153 : std_logic_vector(0 to 0) := (others => '0');
    variable r151 : std_logic_vector(0 to 0) := (others => '0');
    variable r149 : std_logic_vector(0 to 7) := (others => '0');
    variable r147 : std_logic_vector(0 to 0) := (others => '0');
    variable r145 : std_logic_vector(0 to 0) := (others => '0');
    variable r143 : std_logic_vector(0 to 0) := (others => '0');
    variable r141 : std_logic_vector(0 to 0) := (others => '0');
    variable r139 : std_logic_vector(0 to 0) := (others => '0');
    variable r137 : std_logic_vector(0 to 0) := (others => '0');
    variable r135 : std_logic_vector(0 to 0) := (others => '0');
    variable r133 : std_logic_vector(0 to 0) := (others => '0');
    variable r131 : std_logic_vector(0 to 7) := (others => '0');
    variable r129 : std_logic_vector(0 to 0) := (others => '0');
    variable r127 : std_logic_vector(0 to 0) := (others => '0');
    variable r125 : std_logic_vector(0 to 0) := (others => '0');
    variable r123 : std_logic_vector(0 to 0) := (others => '0');
    variable r121 : std_logic_vector(0 to 0) := (others => '0');
    variable r119 : std_logic_vector(0 to 0) := (others => '0');
    variable r117 : std_logic_vector(0 to 0) := (others => '0');
    variable r115 : std_logic_vector(0 to 0) := (others => '0');
    variable r113 : std_logic_vector(0 to 7) := (others => '0');
    variable r111 : std_logic_vector(0 to 0) := (others => '0');
    variable r109 : std_logic_vector(0 to 0) := (others => '0');
    variable r107 : std_logic_vector(0 to 0) := (others => '0');
    variable r105 : std_logic_vector(0 to 0) := (others => '0');
    variable r103 : std_logic_vector(0 to 0) := (others => '0');
    variable r101 : std_logic_vector(0 to 0) := (others => '0');
    variable r99 : std_logic_vector(0 to 0) := (others => '0');
    variable r97 : std_logic_vector(0 to 0) := (others => '0');
    variable r95 : std_logic_vector(0 to 7) := (others => '0');
    variable r93 : std_logic_vector(0 to 0) := (others => '0');
    variable r91 : std_logic_vector(0 to 0) := (others => '0');
    variable r89 : std_logic_vector(0 to 0) := (others => '0');
    variable r87 : std_logic_vector(0 to 0) := (others => '0');
    variable r85 : std_logic_vector(0 to 0) := (others => '0');
    variable r83 : std_logic_vector(0 to 0) := (others => '0');
    variable r81 : std_logic_vector(0 to 0) := (others => '0');
    variable r79 : std_logic_vector(0 to 0) := (others => '0');
    variable r77 : std_logic_vector(0 to 7) := (others => '0');
    variable r75 : std_logic_vector(0 to 0) := (others => '0');
    variable r73 : std_logic_vector(0 to 0) := (others => '0');
    variable r71 : std_logic_vector(0 to 0) := (others => '0');
    variable r69 : std_logic_vector(0 to 0) := (others => '0');
    variable r67 : std_logic_vector(0 to 0) := (others => '0');
    variable r65 : std_logic_vector(0 to 0) := (others => '0');
    variable r63 : std_logic_vector(0 to 0) := (others => '0');
    variable r61 : std_logic_vector(0 to 0) := (others => '0');
    variable r59 : std_logic_vector(0 to 7) := (others => '0');
    variable r57 : std_logic_vector(0 to 0) := (others => '0');
    variable r55 : std_logic_vector(0 to 0) := (others => '0');
    variable r53 : std_logic_vector(0 to 0) := (others => '0');
    variable r51 : std_logic_vector(0 to 0) := (others => '0');
    variable r49 : std_logic_vector(0 to 0) := (others => '0');
    variable r47 : std_logic_vector(0 to 0) := (others => '0');
    variable r45 : std_logic_vector(0 to 0) := (others => '0');
    variable r43 : std_logic_vector(0 to 0) := (others => '0');
    variable r41 : std_logic_vector(0 to 7) := (others => '0');
    variable r39 : std_logic_vector(0 to 0) := (others => '0');
    variable r37 : std_logic_vector(0 to 0) := (others => '0');
    variable r35 : std_logic_vector(0 to 0) := (others => '0');
    variable r33 : std_logic_vector(0 to 0) := (others => '0');
    variable r31 : std_logic_vector(0 to 0) := (others => '0');
    variable r29 : std_logic_vector(0 to 0) := (others => '0');
    variable r27 : std_logic_vector(0 to 0) := (others => '0');
    variable r25 : std_logic_vector(0 to 0) := (others => '0');
    variable r23 : std_logic_vector(0 to 7) := (others => '0');
    variable r21 : std_logic_vector(0 to 0) := (others => '0');
    variable r19 : std_logic_vector(0 to 0) := (others => '0');
    variable r17 : std_logic_vector(0 to 0) := (others => '0');
    variable r15 : std_logic_vector(0 to 0) := (others => '0');
    variable r13 : std_logic_vector(0 to 0) := (others => '0');
    variable r11 : std_logic_vector(0 to 0) := (others => '0');
    variable r9 : std_logic_vector(0 to 0) := (others => '0');
    variable r7 : std_logic_vector(0 to 0) := (others => '0');
    variable EMPTY : std_logic_vector(0 to -1) := (others => '0');
  begin
    r7 := "0";
    r9 := "0";
    r11 := "0";
    r13 := "0";
    r15 := "0";
    r17 := "0";
    r19 := "0";
    r21 := "0";
    r23 := (r7 & r9 & r11 & r13 & r15 & r17 & r19 & r21);
    r25 := "0";
    r27 := "0";
    r29 := "0";
    r31 := "0";
    r33 := "0";
    r35 := "0";
    r37 := "0";
    r39 := "0";
    r41 := (r25 & r27 & r29 & r31 & r33 & r35 & r37 & r39);
    r43 := "0";
    r45 := "0";
    r47 := "0";
    r49 := "0";
    r51 := "0";
    r53 := "0";
    r55 := "0";
    r57 := "0";
    r59 := (r43 & r45 & r47 & r49 & r51 & r53 & r55 & r57);
    r61 := "0";
    r63 := "0";
    r65 := "0";
    r67 := "0";
    r69 := "0";
    r71 := "0";
    r73 := "0";
    r75 := "0";
    r77 := (r61 & r63 & r65 & r67 & r69 & r71 & r73 & r75);
    r79 := "0";
    r81 := "0";
    r83 := "0";
    r85 := "0";
    r87 := "0";
    r89 := "0";
    r91 := "0";
    r93 := "0";
    r95 := (r79 & r81 & r83 & r85 & r87 & r89 & r91 & r93);
    r97 := "0";
    r99 := "0";
    r101 := "0";
    r103 := "0";
    r105 := "0";
    r107 := "0";
    r109 := "0";
    r111 := "0";
    r113 := (r97 & r99 & r101 & r103 & r105 & r107 & r109 & r111);
    r115 := "0";
    r117 := "0";
    r119 := "0";
    r121 := "0";
    r123 := "0";
    r125 := "0";
    r127 := "0";
    r129 := "0";
    r131 := (r115 & r117 & r119 & r121 & r123 & r125 & r127 & r129);
    r133 := "0";
    r135 := "0";
    r137 := "0";
    r139 := "0";
    r141 := "0";
    r143 := "0";
    r145 := "0";
    r147 := "0";
    r149 := (r133 & r135 & r137 & r139 & r141 & r143 & r145 & r147);
    r151 := "0";
    r153 := "0";
    r155 := "0";
    r157 := "0";
    r159 := "0";
    r161 := "0";
    r163 := "0";
    r165 := "0";
    r167 := (r151 & r153 & r155 & r157 & r159 & r161 & r163 & r165);
    r169 := "0";
    r171 := "0";
    r173 := "0";
    r175 := "0";
    r177 := "0";
    r179 := "0";
    r181 := "0";
    r183 := "0";
    r185 := (r169 & r171 & r173 & r175 & r177 & r179 & r181 & r183);
    r187 := "0";
    r189 := "0";
    r191 := "0";
    r193 := "0";
    r195 := "0";
    r197 := "0";
    r199 := "0";
    r201 := "0";
    r203 := (r187 & r189 & r191 & r193 & r195 & r197 & r199 & r201);
    r205 := "0";
    r207 := "0";
    r209 := "0";
    r211 := "0";
    r213 := "0";
    r215 := "0";
    r217 := "0";
    r219 := "0";
    r221 := (r205 & r207 & r209 & r211 & r213 & r215 & r217 & r219);
    r223 := "0";
    r225 := "0";
    r227 := "0";
    r229 := "0";
    r231 := "0";
    r233 := "0";
    r235 := "0";
    r237 := "0";
    r239 := (r223 & r225 & r227 & r229 & r231 & r233 & r235 & r237);
    r241 := "0";
    r243 := "0";
    r245 := "0";
    r247 := "0";
    r249 := "0";
    r251 := "0";
    r253 := "0";
    r255 := "0";
    r257 := (r241 & r243 & r245 & r247 & r249 & r251 & r253 & r255);
    r259 := "0";
    r261 := "0";
    r263 := "0";
    r265 := "0";
    r267 := "0";
    r269 := "0";
    r271 := "0";
    r273 := "0";
    r275 := (r259 & r261 & r263 & r265 & r267 & r269 & r271 & r273);
    r277 := "0";
    r279 := "0";
    r281 := "0";
    r283 := "0";
    r285 := "0";
    r287 := "0";
    r289 := "0";
    r291 := "0";
    r293 := (r277 & r279 & r281 & r283 & r285 & r287 & r289 & r291);
    r295 := "0";
    r297 := "0";
    r299 := "0";
    r301 := "0";
    r303 := "0";
    r305 := "0";
    r307 := "0";
    r309 := "0";
    r311 := (r295 & r297 & r299 & r301 & r303 & r305 & r307 & r309);
    r313 := "0";
    r315 := "0";
    r317 := "0";
    r319 := "0";
    r321 := "0";
    r323 := "0";
    r325 := "0";
    r327 := "0";
    r329 := (r313 & r315 & r317 & r319 & r321 & r323 & r325 & r327);
    r331 := "0";
    r333 := "0";
    r335 := "0";
    r337 := "0";
    r339 := "0";
    r341 := "0";
    r343 := "0";
    r345 := "0";
    r347 := (r331 & r333 & r335 & r337 & r339 & r341 & r343 & r345);
    r349 := "0";
    r351 := "0";
    r353 := "0";
    r355 := "0";
    r357 := "0";
    r359 := "0";
    r361 := "0";
    r363 := "0";
    r365 := (r349 & r351 & r353 & r355 & r357 & r359 & r361 & r363);
    r367 := "0";
    r369 := "0";
    r371 := "0";
    r373 := "0";
    r375 := "0";
    r377 := "0";
    r379 := "0";
    r381 := "0";
    r383 := (r367 & r369 & r371 & r373 & r375 & r377 & r379 & r381);
    r385 := "0";
    r387 := "0";
    r389 := "0";
    r391 := "0";
    r393 := "0";
    r395 := "0";
    r397 := "0";
    r399 := "0";
    r401 := (r385 & r387 & r389 & r391 & r393 & r395 & r397 & r399);
    r403 := "0";
    r405 := "0";
    r407 := "0";
    r409 := "0";
    r411 := "0";
    r413 := "0";
    r415 := "0";
    r417 := "0";
    r419 := (r403 & r405 & r407 & r409 & r411 & r413 & r415 & r417);
    r421 := "0";
    r423 := "0";
    r425 := "0";
    r427 := "0";
    r429 := "0";
    r431 := "0";
    r433 := "0";
    r435 := "0";
    r437 := (r421 & r423 & r425 & r427 & r429 & r431 & r433 & r435);
    r439 := "0";
    r441 := "0";
    r443 := "0";
    r445 := "0";
    r447 := "0";
    r449 := "0";
    r451 := "0";
    r453 := "0";
    r455 := (r439 & r441 & r443 & r445 & r447 & r449 & r451 & r453);
    r457 := "0";
    r459 := "0";
    r461 := "0";
    r463 := "0";
    r465 := "0";
    r467 := "0";
    r469 := "0";
    r471 := "0";
    r473 := (r457 & r459 & r461 & r463 & r465 & r467 & r469 & r471);
    r475 := "0";
    r477 := "0";
    r479 := "0";
    r481 := "0";
    r483 := "0";
    r485 := "0";
    r487 := "0";
    r489 := "0";
    r491 := (r475 & r477 & r479 & r481 & r483 & r485 & r487 & r489);
    r493 := "0";
    r495 := "0";
    r497 := "0";
    r499 := "0";
    r501 := "0";
    r503 := "0";
    r505 := "0";
    r507 := "0";
    r509 := (r493 & r495 & r497 & r499 & r501 & r503 & r505 & r507);
    r511 := "0";
    r513 := "0";
    r515 := "0";
    r517 := "0";
    r519 := "0";
    r521 := "0";
    r523 := "0";
    r525 := "0";
    r527 := (r511 & r513 & r515 & r517 & r519 & r521 & r523 & r525);
    r529 := "0";
    r531 := "0";
    r533 := "0";
    r535 := "0";
    r537 := "0";
    r539 := "0";
    r541 := "0";
    r543 := "0";
    r545 := (r529 & r531 & r533 & r535 & r537 & r539 & r541 & r543);
    r547 := "0";
    r549 := "0";
    r551 := "0";
    r553 := "0";
    r555 := "0";
    r557 := "0";
    r559 := "0";
    r561 := "0";
    r563 := (r547 & r549 & r551 & r553 & r555 & r557 & r559 & r561);
    r565 := "0";
    r567 := "0";
    r569 := "0";
    r571 := "0";
    r573 := "0";
    r575 := "0";
    r577 := "0";
    r579 := "0";
    r581 := (r565 & r567 & r569 & r571 & r573 & r575 & r577 & r579);
    r583 := "0";
    r585 := "0";
    r587 := "0";
    r589 := "0";
    r591 := "0";
    r593 := "0";
    r595 := "0";
    r597 := "0";
    r599 := (r583 & r585 & r587 & r589 & r591 & r593 & r595 & r597);
    r601 := "0";
    r603 := "0";
    r605 := "0";
    r607 := "0";
    r609 := "0";
    r611 := "0";
    r613 := "0";
    r615 := "0";
    r617 := (r601 & r603 & r605 & r607 & r609 & r611 & r613 & r615);
    r619 := "0";
    r621 := "0";
    r623 := "0";
    r625 := "0";
    r627 := "0";
    r629 := "0";
    r631 := "0";
    r633 := "0";
    r635 := (r619 & r621 & r623 & r625 & r627 & r629 & r631 & r633);
    r637 := "0";
    r639 := "0";
    r641 := "0";
    r643 := "0";
    r645 := "0";
    r647 := "0";
    r649 := "0";
    r651 := "0";
    r653 := (r637 & r639 & r641 & r643 & r645 & r647 & r649 & r651);
    r655 := "0";
    r657 := "0";
    r659 := "0";
    r661 := "0";
    r663 := "0";
    r665 := "0";
    r667 := "0";
    r669 := "0";
    r671 := (r655 & r657 & r659 & r661 & r663 & r665 & r667 & r669);
    r673 := "0";
    r675 := "0";
    r677 := "0";
    r679 := "0";
    r681 := "0";
    r683 := "0";
    r685 := "0";
    r687 := "0";
    r689 := (r673 & r675 & r677 & r679 & r681 & r683 & r685 & r687);
    r691 := "0";
    r693 := "0";
    r695 := "0";
    r697 := "0";
    r699 := "0";
    r701 := "0";
    r703 := "0";
    r705 := "0";
    r707 := (r691 & r693 & r695 & r697 & r699 & r701 & r703 & r705);
    r709 := "0";
    r711 := "0";
    r713 := "0";
    r715 := "0";
    r717 := "0";
    r719 := "0";
    r721 := "0";
    r723 := "0";
    r725 := (r709 & r711 & r713 & r715 & r717 & r719 & r721 & r723);
    r727 := "0";
    r729 := "0";
    r731 := "0";
    r733 := "0";
    r735 := "0";
    r737 := "0";
    r739 := "0";
    r741 := "0";
    r743 := (r727 & r729 & r731 & r733 & r735 & r737 & r739 & r741);
    r745 := "0";
    r747 := "0";
    r749 := "0";
    r751 := "0";
    r753 := "0";
    r755 := "0";
    r757 := "0";
    r759 := "0";
    r761 := (r745 & r747 & r749 & r751 & r753 & r755 & r757 & r759);
    r763 := "0";
    r765 := "0";
    r767 := "0";
    r769 := "0";
    r771 := "0";
    r773 := "0";
    r775 := "0";
    r777 := "0";
    r779 := (r763 & r765 & r767 & r769 & r771 & r773 & r775 & r777);
    r781 := "0";
    r783 := "0";
    r785 := "0";
    r787 := "0";
    r789 := "0";
    r791 := "0";
    r793 := "0";
    r795 := "0";
    r797 := (r781 & r783 & r785 & r787 & r789 & r791 & r793 & r795);
    r799 := "0";
    r801 := "0";
    r803 := "0";
    r805 := "0";
    r807 := "0";
    r809 := "0";
    r811 := "0";
    r813 := "0";
    r815 := (r799 & r801 & r803 & r805 & r807 & r809 & r811 & r813);
    r817 := "0";
    r819 := "0";
    r821 := "0";
    r823 := "0";
    r825 := "0";
    r827 := "0";
    r829 := "0";
    r831 := "0";
    r833 := (r817 & r819 & r821 & r823 & r825 & r827 & r829 & r831);
    r835 := "0";
    r837 := "0";
    r839 := "0";
    r841 := "0";
    r843 := "0";
    r845 := "0";
    r847 := "0";
    r849 := "0";
    r851 := (r835 & r837 & r839 & r841 & r843 & r845 & r847 & r849);
    r853 := "0";
    r855 := "0";
    r857 := "0";
    r859 := "0";
    r861 := "0";
    r863 := "0";
    r865 := "0";
    r867 := "0";
    r869 := (r853 & r855 & r857 & r859 & r861 & r863 & r865 & r867);
    r871 := "0";
    r873 := "0";
    r875 := "0";
    r877 := "0";
    r879 := "0";
    r881 := "0";
    r883 := "0";
    r885 := "0";
    r887 := (r871 & r873 & r875 & r877 & r879 & r881 & r883 & r885);
    r889 := "0";
    r891 := "0";
    r893 := "0";
    r895 := "0";
    r897 := "0";
    r899 := "0";
    r901 := "0";
    r903 := "0";
    r905 := (r889 & r891 & r893 & r895 & r897 & r899 & r901 & r903);
    r907 := "0";
    r909 := "0";
    r911 := "0";
    r913 := "0";
    r915 := "0";
    r917 := "0";
    r919 := "0";
    r921 := "0";
    r923 := (r907 & r909 & r911 & r913 & r915 & r917 & r919 & r921);
    r925 := "0";
    r927 := "0";
    r929 := "0";
    r931 := "0";
    r933 := "0";
    r935 := "0";
    r937 := "0";
    r939 := "0";
    r941 := (r925 & r927 & r929 & r931 & r933 & r935 & r937 & r939);
    r943 := "0";
    r945 := "0";
    r947 := "0";
    r949 := "0";
    r951 := "0";
    r953 := "0";
    r955 := "0";
    r957 := "0";
    r959 := (r943 & r945 & r947 & r949 & r951 & r953 & r955 & r957);
    r961 := "0";
    r963 := "0";
    r965 := "0";
    r967 := "0";
    r969 := "0";
    r971 := "0";
    r973 := "0";
    r975 := "0";
    r977 := (r961 & r963 & r965 & r967 & r969 & r971 & r973 & r975);
    r979 := "0";
    r981 := "0";
    r983 := "0";
    r985 := "0";
    r987 := "0";
    r989 := "0";
    r991 := "0";
    r993 := "0";
    r995 := (r979 & r981 & r983 & r985 & r987 & r989 & r991 & r993);
    r997 := "0";
    r999 := "0";
    r1001 := "0";
    r1003 := "0";
    r1005 := "0";
    r1007 := "0";
    r1009 := "0";
    r1011 := "0";
    r1013 := (r997 & r999 & r1001 & r1003 & r1005 & r1007 & r1009 & r1011);
    r1015 := "0";
    r1017 := "0";
    r1019 := "0";
    r1021 := "0";
    r1023 := "0";
    r1025 := "0";
    r1027 := "0";
    r1029 := "0";
    r1031 := (r1015 & r1017 & r1019 & r1021 & r1023 & r1025 & r1027 & r1029);
    r1033 := "0";
    r1035 := "0";
    r1037 := "0";
    r1039 := "0";
    r1041 := "0";
    r1043 := "0";
    r1045 := "0";
    r1047 := "0";
    r1049 := (r1033 & r1035 & r1037 & r1039 & r1041 & r1043 & r1045 & r1047);
    r1051 := "0";
    r1053 := "0";
    r1055 := "0";
    r1057 := "0";
    r1059 := "0";
    r1061 := "0";
    r1063 := "0";
    r1065 := "0";
    r1067 := (r1051 & r1053 & r1055 & r1057 & r1059 & r1061 & r1063 & r1065);
    r1069 := "0";
    r1071 := "0";
    r1073 := "0";
    r1075 := "0";
    r1077 := "0";
    r1079 := "0";
    r1081 := "0";
    r1083 := "0";
    r1085 := (r1069 & r1071 & r1073 & r1075 & r1077 & r1079 & r1081 & r1083);
    r1087 := "0";
    r1089 := "0";
    r1091 := "0";
    r1093 := "0";
    r1095 := "0";
    r1097 := "0";
    r1099 := "0";
    r1101 := "0";
    r1103 := (r1087 & r1089 & r1091 & r1093 & r1095 & r1097 & r1099 & r1101);
    r1105 := "0";
    r1107 := "0";
    r1109 := "0";
    r1111 := "0";
    r1113 := "0";
    r1115 := "0";
    r1117 := "0";
    r1119 := "0";
    r1121 := (r1105 & r1107 & r1109 & r1111 & r1113 & r1115 & r1117 & r1119);
    r1123 := "0";
    r1125 := "0";
    r1127 := "0";
    r1129 := "0";
    r1131 := "0";
    r1133 := "0";
    r1135 := "0";
    r1137 := "0";
    r1139 := (r1123 & r1125 & r1127 & r1129 & r1131 & r1133 & r1135 & r1137);
    r1141 := "0";
    r1143 := "0";
    r1145 := "0";
    r1147 := "0";
    r1149 := "0";
    r1151 := "0";
    r1153 := "0";
    r1155 := "0";
    r1157 := (r1141 & r1143 & r1145 & r1147 & r1149 & r1151 & r1153 & r1155);
    r1158 := (r23 & r41 & r59 & r77 & r95 & r113 & r131 & r149 & r167 & r185 & r203 & r221 & r239 & r257 & r275 & r293 & r311 & r329 & r347 & r365 & r383 & r401 & r419 & r437 & r455 & r473 & r491 & r509 & r527 & r545 & r563 & r581 & r599 & r617 & r635 & r653 & r671 & r689 & r707 & r725 & r743 & r761 & r779 & r797 & r815 & r833 & r851 & r869 & r887 & r905 & r923 & r941 & r959 & r977 & r995 & r1013 & r1031 & r1049 & r1067 & r1085 & r1103 & r1121 & r1139 & r1157);
    return r1158;
  end rewire_zerothoutput_3;

begin
  process (clk)
    variable goto_L3536 : boolean := false;
    variable goto_L3530 : boolean := false;
    variable goto_L1163 : boolean := false;
    variable goto_L1165 : boolean := false;
    variable goto_L0 : boolean := false;
    variable goto_L3537 : boolean := false;
    variable r3529 : std_logic_vector(0 to 127) := (others => '0');
    variable r3525 : std_logic_vector(0 to 511) := (others => '0');
    variable r3521 : std_logic_vector(0 to 127) := (others => '0');
    variable r3230 : std_logic_vector(0 to 127) := (others => '0');
    variable r3227 : std_logic_vector(0 to 127) := (others => '0');
    variable r2936 : std_logic_vector(0 to 127) := (others => '0');
    variable r1183 : std_logic_vector(0 to 511) := (others => '0');
    variable r1182 : std_logic_vector(0 to 63) := (others => '0');
    variable r1181 : std_logic_vector(0 to 63) := (others => '0');
    variable r1180 : std_logic_vector(0 to 127) := (others => '0');
    variable r1179 : std_logic_vector(0 to 127) := (others => '0');
    variable b1176 : boolean := false;
    variable b1174 : boolean := false;
    variable r1172 : std_logic_vector(0 to 63) := (others => '0');
    variable r1170 : std_logic_vector(0 to 63) := (others => '0');
    variable r1164 : std_logic_vector(0 to 127) := (others => '0');
    variable r1162 : std_logic_vector(0 to 127) := (others => '0');
    variable r1159 : std_logic_vector(0 to 511) := (others => '0');
    variable r4 : std_logic_vector(0 to 511) := (others => '0');
    variable EMPTY : std_logic_vector(0 to -1) := (others => '0');
    variable state : control_state := STATE0;
  begin
    if clk'event and clk='1' then
      goto_L3536 := false;
      goto_L3530 := false;
      goto_L1163 := false;
      goto_L1165 := false;
      goto_L0 := false;
      goto_L3537 := false;
      null; -- label L3536
      -- ENTER
      goto_L0 := (state = STATE0);
      if (NOT goto_L0) then
        goto_L1163 := (state = STATE1163);
        if (NOT goto_L1163) then
          goto_L3530 := (state = STATE3530);
          null; -- label L3530
          r3529 := input;
          -- got r@IT in r3529
          r1164 := r3529;
          goto_L1165 := true;
        end if;
        goto_L1165 := goto_L1165;
        if (NOT goto_L1165) then
          null; -- label L1163
          r1162 := input;
          -- got r@IU in r1162
          r1164 := r1162;
          goto_L1165 := true;
        end if;
        goto_L1165 := goto_L1165;
        null; -- label L1165
        -- step in
        -- got x@IP in r1164
        -- final pat
        r1170 := r1164(0 to 63);
        r1172 := r1164(64 to 127);
        b1174 := true;
        b1176 := true;
        r3227 := rewire_key1_2935;
        r3521 := rewire_key2_3229;
        -- got b0@IQ in r1170
        -- got b1@IR in r1172
        r3525 := rewire_buildSalsa256_1178(r3227,r3521,r1170,r1172);
        -- got y@IS in r3525
        output <= r3525;
        state := STATE3530;
        goto_L3537 := true;
      end if;
      goto_L3537 := goto_L3537;
      if (NOT goto_L3537) then
        null; -- label L0
        -- START
        -- foo in
        r1159 := rewire_zerothoutput_3;
        output <= r1159;
        state := STATE1163;
        goto_L3537 := true;
      end if;
      goto_L3537 := goto_L3537;
      null; -- label L3537
      -- EXIT
    end if;
  end process;
end behavioral;
library ieee;
use ieee.std_logic_1164.all;
-- Uncomment the following line if VHDL primitives are in use.
use work.prims.all;
entity main is
  Port ( clk : in std_logic ;
         input : in std_logic_vector (0 to 127);
         output : out std_logic_vector (0 to 511));
end main;
architecture structural of main is
begin
  dev : entity work.rwcomp0(behavioral)
    port map (clk,input,output);
    

end structural;
