library ieee;
use ieee.std_logic_1164.all;
-- Uncomment the following line if VHDL primitives are in use.
use work.prims.all;
entity rwcomp0 is
  Port ( clk : in std_logic ;
         input : in std_logic_vector (0 to 9);
         output : out std_logic_vector (0 to 17));
end rwcomp0;

architecture behavioral of rwcomp0 is
  type control_state is (STATE0,STATE182,STATE314,STATE705,STATE814,STATE1189,STATE1506,STATE1723,STATE1927,STATE2135,STATE2339,STATE2547,STATE2676,STATE2862,STATE3048,STATE3234,STATE3408,STATE3517,STATE3628,STATE3737,STATE3848,STATE3943,STATE4004,STATE4091,STATE4285,STATE4422,STATE4521,STATE4703,STATE4885,STATE5026,STATE5128,STATE5383,STATE5427);
  function rewire_csFlag_4235(r4236 : std_logic_vector) return std_logic_vector;
  function rewire_zsFlag_4191(r4192 : std_logic_vector) return std_logic_vector;
  function rewire_pcSave_4147(r4148 : std_logic_vector) return std_logic_vector;
  function rewire_setIackOut_4058(r4059 : std_logic_vector ; r4060 : std_logic_vector) return std_logic_vector;
  function rewire_setR3_1349(r1350 : std_logic_vector ; r1351 : std_logic_vector) return std_logic_vector;
  function rewire_setR2_1306(r1307 : std_logic_vector ; r1308 : std_logic_vector) return std_logic_vector;
  function rewire_setR1_1262(r1263 : std_logic_vector ; r1264 : std_logic_vector) return std_logic_vector;
  function rewire_setR0_1218(r1219 : std_logic_vector ; r1220 : std_logic_vector) return std_logic_vector;
  function rewire_setPC_1124(r1125 : std_logic_vector ; r1126 : std_logic_vector) return std_logic_vector;
  function rewire_setDataOut_1090(r1091 : std_logic_vector ; r1092 : std_logic_vector) return std_logic_vector;
  function rewire_r3_1046(r1047 : std_logic_vector) return std_logic_vector;
  function rewire_r2_1008(r1009 : std_logic_vector) return std_logic_vector;
  function rewire_r1_969(r970 : std_logic_vector) return std_logic_vector;
  function rewire_r0_930(r931 : std_logic_vector) return std_logic_vector;
  function rewire_mkReg_883(r884 : std_logic_vector ; r885 : std_logic_vector) return std_logic_vector;
  function rewire_setWeOut_853(r854 : std_logic_vector ; r855 : std_logic_vector) return std_logic_vector;
  function rewire_setAddrOut_782(r783 : std_logic_vector ; r784 : std_logic_vector) return std_logic_vector;
  function rewire_dataIn_717(r718 : std_logic_vector) return std_logic_vector;
  function rewire_setCSave_657(r658 : std_logic_vector ; r659 : std_logic_vector) return std_logic_vector;
  function rewire_setZSave_615(r616 : std_logic_vector ; r617 : std_logic_vector) return std_logic_vector;
  function rewire_setPCSave_573(r574 : std_logic_vector ; r575 : std_logic_vector) return std_logic_vector;
  function rewire_cFlag_536(r537 : std_logic_vector) return std_logic_vector;
  function rewire_zFlag_499(r500 : std_logic_vector) return std_logic_vector;
  function rewire_pc_462(r463 : std_logic_vector) return std_logic_vector;
  function rewire_setIEFlag_419(r420 : std_logic_vector ; r421 : std_logic_vector) return std_logic_vector;
  function rewire_intIn_387(r388 : std_logic_vector) return std_logic_vector;
  function rewire_rstIn_264(r265 : std_logic_vector) return std_logic_vector;
  function rewire_inputs_229(r230 : std_logic_vector) return std_logic_vector;
  function rewire_setInputs_185(r186 : std_logic_vector ; r187 : std_logic_vector) return std_logic_vector;
  function rewire_outputs_144(r145 : std_logic_vector) return std_logic_vector;
  function rewire_initOutputs_127 return std_logic_vector;
  function rewire_setOutputs_91(r92 : std_logic_vector ; r93 : std_logic_vector) return std_logic_vector;
  function rewire_setZFlag_48(r49 : std_logic_vector ; r50 : std_logic_vector) return std_logic_vector;
  function rewire_setCFlag_5(r6 : std_logic_vector ; r7 : std_logic_vector) return std_logic_vector;

  function rewire_csFlag_4235(r4236 : std_logic_vector) return std_logic_vector
  is
    variable b4266 : boolean := false;
    variable b4265 : boolean := false;
    variable b4264 : boolean := false;
    variable b4263 : boolean := false;
    variable b4262 : boolean := false;
    variable b4261 : boolean := false;
    variable b4260 : boolean := false;
    variable b4259 : boolean := false;
    variable b4258 : boolean := false;
    variable b4257 : boolean := false;
    variable b4256 : boolean := false;
    variable b4255 : boolean := false;
    variable b4254 : boolean := false;
    variable b4253 : boolean := false;
    variable r4252 : std_logic_vector(0 to 7) := (others => '0');
    variable r4251 : std_logic_vector(0 to 7) := (others => '0');
    variable r4250 : std_logic_vector(0 to 7) := (others => '0');
    variable r4249 : std_logic_vector(0 to 7) := (others => '0');
    variable r4248 : std_logic_vector(0 to 7) := (others => '0');
    variable r4247 : std_logic_vector(0 to 0) := (others => '0');
    variable r4246 : std_logic_vector(0 to 0) := (others => '0');
    variable r4245 : std_logic_vector(0 to 7) := (others => '0');
    variable r4244 : std_logic_vector(0 to 0) := (others => '0');
    variable r4243 : std_logic_vector(0 to 0) := (others => '0');
    variable r4242 : std_logic_vector(0 to 0) := (others => '0');
    variable r4241 : std_logic_vector(0 to 17) := (others => '0');
    variable r4240 : std_logic_vector(0 to 9) := (others => '0');
    variable b4239 : boolean := false;
    variable r4238 : std_logic_vector(0 to 0) := (others => '0');
  begin
    null;
    b4239 := true;
    r4240 := r4236(0 to 9);
    r4241 := r4236(10 to 27);
    r4242 := r4236(28 to 28);
    r4243 := r4236(29 to 29);
    r4244 := r4236(30 to 30);
    r4245 := r4236(31 to 38);
    r4246 := r4236(39 to 39);
    r4247 := r4236(40 to 40);
    r4248 := r4236(41 to 48);
    r4249 := r4236(49 to 56);
    r4250 := r4236(57 to 64);
    r4251 := r4236(65 to 72);
    r4252 := r4236(73 to 80);
    b4253 := true;
    b4254 := true;
    b4255 := true;
    b4256 := true;
    b4257 := true;
    b4258 := true;
    b4259 := true;
    b4260 := true;
    b4261 := true;
    b4262 := true;
    b4263 := true;
    b4264 := true;
    b4265 := true;
    b4266 := (b4253 AND (b4254 AND (b4255 AND (b4256 AND (b4257 AND (b4258 AND (b4259 AND (b4260 AND (b4261 AND (b4262 AND (b4263 AND (b4264 AND b4265))))))))))));
    if b4266 then
      null;
      r4238 := r4247;
    end if;
    return r4238;
  end rewire_csFlag_4235;
  function rewire_zsFlag_4191(r4192 : std_logic_vector) return std_logic_vector
  is
    variable b4222 : boolean := false;
    variable b4221 : boolean := false;
    variable b4220 : boolean := false;
    variable b4219 : boolean := false;
    variable b4218 : boolean := false;
    variable b4217 : boolean := false;
    variable b4216 : boolean := false;
    variable b4215 : boolean := false;
    variable b4214 : boolean := false;
    variable b4213 : boolean := false;
    variable b4212 : boolean := false;
    variable b4211 : boolean := false;
    variable b4210 : boolean := false;
    variable b4209 : boolean := false;
    variable r4208 : std_logic_vector(0 to 7) := (others => '0');
    variable r4207 : std_logic_vector(0 to 7) := (others => '0');
    variable r4206 : std_logic_vector(0 to 7) := (others => '0');
    variable r4205 : std_logic_vector(0 to 7) := (others => '0');
    variable r4204 : std_logic_vector(0 to 7) := (others => '0');
    variable r4203 : std_logic_vector(0 to 0) := (others => '0');
    variable r4202 : std_logic_vector(0 to 0) := (others => '0');
    variable r4201 : std_logic_vector(0 to 7) := (others => '0');
    variable r4200 : std_logic_vector(0 to 0) := (others => '0');
    variable r4199 : std_logic_vector(0 to 0) := (others => '0');
    variable r4198 : std_logic_vector(0 to 0) := (others => '0');
    variable r4197 : std_logic_vector(0 to 17) := (others => '0');
    variable r4196 : std_logic_vector(0 to 9) := (others => '0');
    variable b4195 : boolean := false;
    variable r4194 : std_logic_vector(0 to 0) := (others => '0');
  begin
    null;
    b4195 := true;
    r4196 := r4192(0 to 9);
    r4197 := r4192(10 to 27);
    r4198 := r4192(28 to 28);
    r4199 := r4192(29 to 29);
    r4200 := r4192(30 to 30);
    r4201 := r4192(31 to 38);
    r4202 := r4192(39 to 39);
    r4203 := r4192(40 to 40);
    r4204 := r4192(41 to 48);
    r4205 := r4192(49 to 56);
    r4206 := r4192(57 to 64);
    r4207 := r4192(65 to 72);
    r4208 := r4192(73 to 80);
    b4209 := true;
    b4210 := true;
    b4211 := true;
    b4212 := true;
    b4213 := true;
    b4214 := true;
    b4215 := true;
    b4216 := true;
    b4217 := true;
    b4218 := true;
    b4219 := true;
    b4220 := true;
    b4221 := true;
    b4222 := (b4209 AND (b4210 AND (b4211 AND (b4212 AND (b4213 AND (b4214 AND (b4215 AND (b4216 AND (b4217 AND (b4218 AND (b4219 AND (b4220 AND b4221))))))))))));
    if b4222 then
      null;
      r4194 := r4202;
    end if;
    return r4194;
  end rewire_zsFlag_4191;
  function rewire_pcSave_4147(r4148 : std_logic_vector) return std_logic_vector
  is
    variable b4178 : boolean := false;
    variable b4177 : boolean := false;
    variable b4176 : boolean := false;
    variable b4175 : boolean := false;
    variable b4174 : boolean := false;
    variable b4173 : boolean := false;
    variable b4172 : boolean := false;
    variable b4171 : boolean := false;
    variable b4170 : boolean := false;
    variable b4169 : boolean := false;
    variable b4168 : boolean := false;
    variable b4167 : boolean := false;
    variable b4166 : boolean := false;
    variable b4165 : boolean := false;
    variable r4164 : std_logic_vector(0 to 7) := (others => '0');
    variable r4163 : std_logic_vector(0 to 7) := (others => '0');
    variable r4162 : std_logic_vector(0 to 7) := (others => '0');
    variable r4161 : std_logic_vector(0 to 7) := (others => '0');
    variable r4160 : std_logic_vector(0 to 7) := (others => '0');
    variable r4159 : std_logic_vector(0 to 0) := (others => '0');
    variable r4158 : std_logic_vector(0 to 0) := (others => '0');
    variable r4157 : std_logic_vector(0 to 7) := (others => '0');
    variable r4156 : std_logic_vector(0 to 0) := (others => '0');
    variable r4155 : std_logic_vector(0 to 0) := (others => '0');
    variable r4154 : std_logic_vector(0 to 0) := (others => '0');
    variable r4153 : std_logic_vector(0 to 17) := (others => '0');
    variable r4152 : std_logic_vector(0 to 9) := (others => '0');
    variable b4151 : boolean := false;
    variable r4150 : std_logic_vector(0 to 7) := (others => '0');
  begin
    null;
    b4151 := true;
    r4152 := r4148(0 to 9);
    r4153 := r4148(10 to 27);
    r4154 := r4148(28 to 28);
    r4155 := r4148(29 to 29);
    r4156 := r4148(30 to 30);
    r4157 := r4148(31 to 38);
    r4158 := r4148(39 to 39);
    r4159 := r4148(40 to 40);
    r4160 := r4148(41 to 48);
    r4161 := r4148(49 to 56);
    r4162 := r4148(57 to 64);
    r4163 := r4148(65 to 72);
    r4164 := r4148(73 to 80);
    b4165 := true;
    b4166 := true;
    b4167 := true;
    b4168 := true;
    b4169 := true;
    b4170 := true;
    b4171 := true;
    b4172 := true;
    b4173 := true;
    b4174 := true;
    b4175 := true;
    b4176 := true;
    b4177 := true;
    b4178 := (b4165 AND (b4166 AND (b4167 AND (b4168 AND (b4169 AND (b4170 AND (b4171 AND (b4172 AND (b4173 AND (b4174 AND (b4175 AND (b4176 AND b4177))))))))))));
    if b4178 then
      null;
      r4150 := r4160;
    end if;
    return r4150;
  end rewire_pcSave_4147;
  function rewire_setIackOut_4058(r4059 : std_logic_vector ; r4060 : std_logic_vector) return std_logic_vector
  is
    variable r4074 : std_logic_vector(0 to 17) := (others => '0');
    variable EMPTY : std_logic_vector(0 to -1) := (others => '0');
    variable b4072 : boolean := false;
    variable b4071 : boolean := false;
    variable b4070 : boolean := false;
    variable b4069 : boolean := false;
    variable b4068 : boolean := false;
    variable r4067 : std_logic_vector(0 to 0) := (others => '0');
    variable r4066 : std_logic_vector(0 to 0) := (others => '0');
    variable r4065 : std_logic_vector(0 to 7) := (others => '0');
    variable r4064 : std_logic_vector(0 to 7) := (others => '0');
    variable b4063 : boolean := false;
    variable r4062 : std_logic_vector(0 to 17) := (others => '0');
  begin
    null;
    b4063 := true;
    r4064 := r4059(0 to 7);
    r4065 := r4059(8 to 15);
    r4066 := r4059(16 to 16);
    r4067 := r4059(17 to 17);
    b4068 := true;
    b4069 := true;
    b4070 := true;
    b4071 := true;
    b4072 := (b4068 AND (b4069 AND (b4070 AND b4071)));
    if b4072 then
      null;
      null;
      null;
      null;
      r4074 := (r4064 & r4065 & r4066 & r4060);
      r4062 := r4074;
    end if;
    return r4062;
  end rewire_setIackOut_4058;
  function rewire_setR3_1349(r1350 : std_logic_vector ; r1351 : std_logic_vector) return std_logic_vector
  is
    variable r1383 : std_logic_vector(0 to 80) := (others => '0');
    variable EMPTY : std_logic_vector(0 to -1) := (others => '0');
    variable b1381 : boolean := false;
    variable b1380 : boolean := false;
    variable b1379 : boolean := false;
    variable b1378 : boolean := false;
    variable b1377 : boolean := false;
    variable b1376 : boolean := false;
    variable b1375 : boolean := false;
    variable b1374 : boolean := false;
    variable b1373 : boolean := false;
    variable b1372 : boolean := false;
    variable b1371 : boolean := false;
    variable b1370 : boolean := false;
    variable b1369 : boolean := false;
    variable b1368 : boolean := false;
    variable r1367 : std_logic_vector(0 to 7) := (others => '0');
    variable r1366 : std_logic_vector(0 to 7) := (others => '0');
    variable r1365 : std_logic_vector(0 to 7) := (others => '0');
    variable r1364 : std_logic_vector(0 to 7) := (others => '0');
    variable r1363 : std_logic_vector(0 to 7) := (others => '0');
    variable r1362 : std_logic_vector(0 to 0) := (others => '0');
    variable r1361 : std_logic_vector(0 to 0) := (others => '0');
    variable r1360 : std_logic_vector(0 to 7) := (others => '0');
    variable r1359 : std_logic_vector(0 to 0) := (others => '0');
    variable r1358 : std_logic_vector(0 to 0) := (others => '0');
    variable r1357 : std_logic_vector(0 to 0) := (others => '0');
    variable r1356 : std_logic_vector(0 to 17) := (others => '0');
    variable r1355 : std_logic_vector(0 to 9) := (others => '0');
    variable b1354 : boolean := false;
    variable r1353 : std_logic_vector(0 to 80) := (others => '0');
  begin
    null;
    b1354 := true;
    r1355 := r1350(0 to 9);
    r1356 := r1350(10 to 27);
    r1357 := r1350(28 to 28);
    r1358 := r1350(29 to 29);
    r1359 := r1350(30 to 30);
    r1360 := r1350(31 to 38);
    r1361 := r1350(39 to 39);
    r1362 := r1350(40 to 40);
    r1363 := r1350(41 to 48);
    r1364 := r1350(49 to 56);
    r1365 := r1350(57 to 64);
    r1366 := r1350(65 to 72);
    r1367 := r1350(73 to 80);
    b1368 := true;
    b1369 := true;
    b1370 := true;
    b1371 := true;
    b1372 := true;
    b1373 := true;
    b1374 := true;
    b1375 := true;
    b1376 := true;
    b1377 := true;
    b1378 := true;
    b1379 := true;
    b1380 := true;
    b1381 := (b1368 AND (b1369 AND (b1370 AND (b1371 AND (b1372 AND (b1373 AND (b1374 AND (b1375 AND (b1376 AND (b1377 AND (b1378 AND (b1379 AND b1380))))))))))));
    if b1381 then
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      r1383 := (r1355 & r1356 & r1357 & r1358 & r1359 & r1360 & r1361 & r1362 & r1363 & r1364 & r1365 & r1366 & r1351);
      r1353 := r1383;
    end if;
    return r1353;
  end rewire_setR3_1349;
  function rewire_setR2_1306(r1307 : std_logic_vector ; r1308 : std_logic_vector) return std_logic_vector
  is
    variable r1340 : std_logic_vector(0 to 80) := (others => '0');
    variable EMPTY : std_logic_vector(0 to -1) := (others => '0');
    variable b1338 : boolean := false;
    variable b1337 : boolean := false;
    variable b1336 : boolean := false;
    variable b1335 : boolean := false;
    variable b1334 : boolean := false;
    variable b1333 : boolean := false;
    variable b1332 : boolean := false;
    variable b1331 : boolean := false;
    variable b1330 : boolean := false;
    variable b1329 : boolean := false;
    variable b1328 : boolean := false;
    variable b1327 : boolean := false;
    variable b1326 : boolean := false;
    variable b1325 : boolean := false;
    variable r1324 : std_logic_vector(0 to 7) := (others => '0');
    variable r1323 : std_logic_vector(0 to 7) := (others => '0');
    variable r1322 : std_logic_vector(0 to 7) := (others => '0');
    variable r1321 : std_logic_vector(0 to 7) := (others => '0');
    variable r1320 : std_logic_vector(0 to 7) := (others => '0');
    variable r1319 : std_logic_vector(0 to 0) := (others => '0');
    variable r1318 : std_logic_vector(0 to 0) := (others => '0');
    variable r1317 : std_logic_vector(0 to 7) := (others => '0');
    variable r1316 : std_logic_vector(0 to 0) := (others => '0');
    variable r1315 : std_logic_vector(0 to 0) := (others => '0');
    variable r1314 : std_logic_vector(0 to 0) := (others => '0');
    variable r1313 : std_logic_vector(0 to 17) := (others => '0');
    variable r1312 : std_logic_vector(0 to 9) := (others => '0');
    variable b1311 : boolean := false;
    variable r1310 : std_logic_vector(0 to 80) := (others => '0');
  begin
    null;
    b1311 := true;
    r1312 := r1307(0 to 9);
    r1313 := r1307(10 to 27);
    r1314 := r1307(28 to 28);
    r1315 := r1307(29 to 29);
    r1316 := r1307(30 to 30);
    r1317 := r1307(31 to 38);
    r1318 := r1307(39 to 39);
    r1319 := r1307(40 to 40);
    r1320 := r1307(41 to 48);
    r1321 := r1307(49 to 56);
    r1322 := r1307(57 to 64);
    r1323 := r1307(65 to 72);
    r1324 := r1307(73 to 80);
    b1325 := true;
    b1326 := true;
    b1327 := true;
    b1328 := true;
    b1329 := true;
    b1330 := true;
    b1331 := true;
    b1332 := true;
    b1333 := true;
    b1334 := true;
    b1335 := true;
    b1336 := true;
    b1337 := true;
    b1338 := (b1325 AND (b1326 AND (b1327 AND (b1328 AND (b1329 AND (b1330 AND (b1331 AND (b1332 AND (b1333 AND (b1334 AND (b1335 AND (b1336 AND b1337))))))))))));
    if b1338 then
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      r1340 := (r1312 & r1313 & r1314 & r1315 & r1316 & r1317 & r1318 & r1319 & r1320 & r1321 & r1322 & r1308 & r1324);
      r1310 := r1340;
    end if;
    return r1310;
  end rewire_setR2_1306;
  function rewire_setR1_1262(r1263 : std_logic_vector ; r1264 : std_logic_vector) return std_logic_vector
  is
    variable r1296 : std_logic_vector(0 to 80) := (others => '0');
    variable EMPTY : std_logic_vector(0 to -1) := (others => '0');
    variable b1294 : boolean := false;
    variable b1293 : boolean := false;
    variable b1292 : boolean := false;
    variable b1291 : boolean := false;
    variable b1290 : boolean := false;
    variable b1289 : boolean := false;
    variable b1288 : boolean := false;
    variable b1287 : boolean := false;
    variable b1286 : boolean := false;
    variable b1285 : boolean := false;
    variable b1284 : boolean := false;
    variable b1283 : boolean := false;
    variable b1282 : boolean := false;
    variable b1281 : boolean := false;
    variable r1280 : std_logic_vector(0 to 7) := (others => '0');
    variable r1279 : std_logic_vector(0 to 7) := (others => '0');
    variable r1278 : std_logic_vector(0 to 7) := (others => '0');
    variable r1277 : std_logic_vector(0 to 7) := (others => '0');
    variable r1276 : std_logic_vector(0 to 7) := (others => '0');
    variable r1275 : std_logic_vector(0 to 0) := (others => '0');
    variable r1274 : std_logic_vector(0 to 0) := (others => '0');
    variable r1273 : std_logic_vector(0 to 7) := (others => '0');
    variable r1272 : std_logic_vector(0 to 0) := (others => '0');
    variable r1271 : std_logic_vector(0 to 0) := (others => '0');
    variable r1270 : std_logic_vector(0 to 0) := (others => '0');
    variable r1269 : std_logic_vector(0 to 17) := (others => '0');
    variable r1268 : std_logic_vector(0 to 9) := (others => '0');
    variable b1267 : boolean := false;
    variable r1266 : std_logic_vector(0 to 80) := (others => '0');
  begin
    null;
    b1267 := true;
    r1268 := r1263(0 to 9);
    r1269 := r1263(10 to 27);
    r1270 := r1263(28 to 28);
    r1271 := r1263(29 to 29);
    r1272 := r1263(30 to 30);
    r1273 := r1263(31 to 38);
    r1274 := r1263(39 to 39);
    r1275 := r1263(40 to 40);
    r1276 := r1263(41 to 48);
    r1277 := r1263(49 to 56);
    r1278 := r1263(57 to 64);
    r1279 := r1263(65 to 72);
    r1280 := r1263(73 to 80);
    b1281 := true;
    b1282 := true;
    b1283 := true;
    b1284 := true;
    b1285 := true;
    b1286 := true;
    b1287 := true;
    b1288 := true;
    b1289 := true;
    b1290 := true;
    b1291 := true;
    b1292 := true;
    b1293 := true;
    b1294 := (b1281 AND (b1282 AND (b1283 AND (b1284 AND (b1285 AND (b1286 AND (b1287 AND (b1288 AND (b1289 AND (b1290 AND (b1291 AND (b1292 AND b1293))))))))))));
    if b1294 then
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      r1296 := (r1268 & r1269 & r1270 & r1271 & r1272 & r1273 & r1274 & r1275 & r1276 & r1277 & r1264 & r1279 & r1280);
      r1266 := r1296;
    end if;
    return r1266;
  end rewire_setR1_1262;
  function rewire_setR0_1218(r1219 : std_logic_vector ; r1220 : std_logic_vector) return std_logic_vector
  is
    variable r1252 : std_logic_vector(0 to 80) := (others => '0');
    variable EMPTY : std_logic_vector(0 to -1) := (others => '0');
    variable b1250 : boolean := false;
    variable b1249 : boolean := false;
    variable b1248 : boolean := false;
    variable b1247 : boolean := false;
    variable b1246 : boolean := false;
    variable b1245 : boolean := false;
    variable b1244 : boolean := false;
    variable b1243 : boolean := false;
    variable b1242 : boolean := false;
    variable b1241 : boolean := false;
    variable b1240 : boolean := false;
    variable b1239 : boolean := false;
    variable b1238 : boolean := false;
    variable b1237 : boolean := false;
    variable r1236 : std_logic_vector(0 to 7) := (others => '0');
    variable r1235 : std_logic_vector(0 to 7) := (others => '0');
    variable r1234 : std_logic_vector(0 to 7) := (others => '0');
    variable r1233 : std_logic_vector(0 to 7) := (others => '0');
    variable r1232 : std_logic_vector(0 to 7) := (others => '0');
    variable r1231 : std_logic_vector(0 to 0) := (others => '0');
    variable r1230 : std_logic_vector(0 to 0) := (others => '0');
    variable r1229 : std_logic_vector(0 to 7) := (others => '0');
    variable r1228 : std_logic_vector(0 to 0) := (others => '0');
    variable r1227 : std_logic_vector(0 to 0) := (others => '0');
    variable r1226 : std_logic_vector(0 to 0) := (others => '0');
    variable r1225 : std_logic_vector(0 to 17) := (others => '0');
    variable r1224 : std_logic_vector(0 to 9) := (others => '0');
    variable b1223 : boolean := false;
    variable r1222 : std_logic_vector(0 to 80) := (others => '0');
  begin
    null;
    b1223 := true;
    r1224 := r1219(0 to 9);
    r1225 := r1219(10 to 27);
    r1226 := r1219(28 to 28);
    r1227 := r1219(29 to 29);
    r1228 := r1219(30 to 30);
    r1229 := r1219(31 to 38);
    r1230 := r1219(39 to 39);
    r1231 := r1219(40 to 40);
    r1232 := r1219(41 to 48);
    r1233 := r1219(49 to 56);
    r1234 := r1219(57 to 64);
    r1235 := r1219(65 to 72);
    r1236 := r1219(73 to 80);
    b1237 := true;
    b1238 := true;
    b1239 := true;
    b1240 := true;
    b1241 := true;
    b1242 := true;
    b1243 := true;
    b1244 := true;
    b1245 := true;
    b1246 := true;
    b1247 := true;
    b1248 := true;
    b1249 := true;
    b1250 := (b1237 AND (b1238 AND (b1239 AND (b1240 AND (b1241 AND (b1242 AND (b1243 AND (b1244 AND (b1245 AND (b1246 AND (b1247 AND (b1248 AND b1249))))))))))));
    if b1250 then
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      r1252 := (r1224 & r1225 & r1226 & r1227 & r1228 & r1229 & r1230 & r1231 & r1232 & r1220 & r1234 & r1235 & r1236);
      r1222 := r1252;
    end if;
    return r1222;
  end rewire_setR0_1218;
  function rewire_setPC_1124(r1125 : std_logic_vector ; r1126 : std_logic_vector) return std_logic_vector
  is
    variable r1158 : std_logic_vector(0 to 80) := (others => '0');
    variable EMPTY : std_logic_vector(0 to -1) := (others => '0');
    variable b1156 : boolean := false;
    variable b1155 : boolean := false;
    variable b1154 : boolean := false;
    variable b1153 : boolean := false;
    variable b1152 : boolean := false;
    variable b1151 : boolean := false;
    variable b1150 : boolean := false;
    variable b1149 : boolean := false;
    variable b1148 : boolean := false;
    variable b1147 : boolean := false;
    variable b1146 : boolean := false;
    variable b1145 : boolean := false;
    variable b1144 : boolean := false;
    variable b1143 : boolean := false;
    variable r1142 : std_logic_vector(0 to 7) := (others => '0');
    variable r1141 : std_logic_vector(0 to 7) := (others => '0');
    variable r1140 : std_logic_vector(0 to 7) := (others => '0');
    variable r1139 : std_logic_vector(0 to 7) := (others => '0');
    variable r1138 : std_logic_vector(0 to 7) := (others => '0');
    variable r1137 : std_logic_vector(0 to 0) := (others => '0');
    variable r1136 : std_logic_vector(0 to 0) := (others => '0');
    variable r1135 : std_logic_vector(0 to 7) := (others => '0');
    variable r1134 : std_logic_vector(0 to 0) := (others => '0');
    variable r1133 : std_logic_vector(0 to 0) := (others => '0');
    variable r1132 : std_logic_vector(0 to 0) := (others => '0');
    variable r1131 : std_logic_vector(0 to 17) := (others => '0');
    variable r1130 : std_logic_vector(0 to 9) := (others => '0');
    variable b1129 : boolean := false;
    variable r1128 : std_logic_vector(0 to 80) := (others => '0');
  begin
    null;
    b1129 := true;
    r1130 := r1125(0 to 9);
    r1131 := r1125(10 to 27);
    r1132 := r1125(28 to 28);
    r1133 := r1125(29 to 29);
    r1134 := r1125(30 to 30);
    r1135 := r1125(31 to 38);
    r1136 := r1125(39 to 39);
    r1137 := r1125(40 to 40);
    r1138 := r1125(41 to 48);
    r1139 := r1125(49 to 56);
    r1140 := r1125(57 to 64);
    r1141 := r1125(65 to 72);
    r1142 := r1125(73 to 80);
    b1143 := true;
    b1144 := true;
    b1145 := true;
    b1146 := true;
    b1147 := true;
    b1148 := true;
    b1149 := true;
    b1150 := true;
    b1151 := true;
    b1152 := true;
    b1153 := true;
    b1154 := true;
    b1155 := true;
    b1156 := (b1143 AND (b1144 AND (b1145 AND (b1146 AND (b1147 AND (b1148 AND (b1149 AND (b1150 AND (b1151 AND (b1152 AND (b1153 AND (b1154 AND b1155))))))))))));
    if b1156 then
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      r1158 := (r1130 & r1131 & r1132 & r1133 & r1134 & r1126 & r1136 & r1137 & r1138 & r1139 & r1140 & r1141 & r1142);
      r1128 := r1158;
    end if;
    return r1128;
  end rewire_setPC_1124;
  function rewire_setDataOut_1090(r1091 : std_logic_vector ; r1092 : std_logic_vector) return std_logic_vector
  is
    variable r1106 : std_logic_vector(0 to 17) := (others => '0');
    variable EMPTY : std_logic_vector(0 to -1) := (others => '0');
    variable b1104 : boolean := false;
    variable b1103 : boolean := false;
    variable b1102 : boolean := false;
    variable b1101 : boolean := false;
    variable b1100 : boolean := false;
    variable r1099 : std_logic_vector(0 to 0) := (others => '0');
    variable r1098 : std_logic_vector(0 to 0) := (others => '0');
    variable r1097 : std_logic_vector(0 to 7) := (others => '0');
    variable r1096 : std_logic_vector(0 to 7) := (others => '0');
    variable b1095 : boolean := false;
    variable r1094 : std_logic_vector(0 to 17) := (others => '0');
  begin
    null;
    b1095 := true;
    r1096 := r1091(0 to 7);
    r1097 := r1091(8 to 15);
    r1098 := r1091(16 to 16);
    r1099 := r1091(17 to 17);
    b1100 := true;
    b1101 := true;
    b1102 := true;
    b1103 := true;
    b1104 := (b1100 AND (b1101 AND (b1102 AND b1103)));
    if b1104 then
      null;
      null;
      null;
      null;
      r1106 := (r1096 & r1092 & r1098 & r1099);
      r1094 := r1106;
    end if;
    return r1094;
  end rewire_setDataOut_1090;
  function rewire_r3_1046(r1047 : std_logic_vector) return std_logic_vector
  is
    variable b1077 : boolean := false;
    variable b1076 : boolean := false;
    variable b1075 : boolean := false;
    variable b1074 : boolean := false;
    variable b1073 : boolean := false;
    variable b1072 : boolean := false;
    variable b1071 : boolean := false;
    variable b1070 : boolean := false;
    variable b1069 : boolean := false;
    variable b1068 : boolean := false;
    variable b1067 : boolean := false;
    variable b1066 : boolean := false;
    variable b1065 : boolean := false;
    variable b1064 : boolean := false;
    variable r1063 : std_logic_vector(0 to 7) := (others => '0');
    variable r1062 : std_logic_vector(0 to 7) := (others => '0');
    variable r1061 : std_logic_vector(0 to 7) := (others => '0');
    variable r1060 : std_logic_vector(0 to 7) := (others => '0');
    variable r1059 : std_logic_vector(0 to 7) := (others => '0');
    variable r1058 : std_logic_vector(0 to 0) := (others => '0');
    variable r1057 : std_logic_vector(0 to 0) := (others => '0');
    variable r1056 : std_logic_vector(0 to 7) := (others => '0');
    variable r1055 : std_logic_vector(0 to 0) := (others => '0');
    variable r1054 : std_logic_vector(0 to 0) := (others => '0');
    variable r1053 : std_logic_vector(0 to 0) := (others => '0');
    variable r1052 : std_logic_vector(0 to 17) := (others => '0');
    variable r1051 : std_logic_vector(0 to 9) := (others => '0');
    variable b1050 : boolean := false;
    variable r1049 : std_logic_vector(0 to 7) := (others => '0');
  begin
    null;
    b1050 := true;
    r1051 := r1047(0 to 9);
    r1052 := r1047(10 to 27);
    r1053 := r1047(28 to 28);
    r1054 := r1047(29 to 29);
    r1055 := r1047(30 to 30);
    r1056 := r1047(31 to 38);
    r1057 := r1047(39 to 39);
    r1058 := r1047(40 to 40);
    r1059 := r1047(41 to 48);
    r1060 := r1047(49 to 56);
    r1061 := r1047(57 to 64);
    r1062 := r1047(65 to 72);
    r1063 := r1047(73 to 80);
    b1064 := true;
    b1065 := true;
    b1066 := true;
    b1067 := true;
    b1068 := true;
    b1069 := true;
    b1070 := true;
    b1071 := true;
    b1072 := true;
    b1073 := true;
    b1074 := true;
    b1075 := true;
    b1076 := true;
    b1077 := (b1064 AND (b1065 AND (b1066 AND (b1067 AND (b1068 AND (b1069 AND (b1070 AND (b1071 AND (b1072 AND (b1073 AND (b1074 AND (b1075 AND b1076))))))))))));
    if b1077 then
      null;
      r1049 := r1063;
    end if;
    return r1049;
  end rewire_r3_1046;
  function rewire_r2_1008(r1009 : std_logic_vector) return std_logic_vector
  is
    variable b1039 : boolean := false;
    variable b1038 : boolean := false;
    variable b1037 : boolean := false;
    variable b1036 : boolean := false;
    variable b1035 : boolean := false;
    variable b1034 : boolean := false;
    variable b1033 : boolean := false;
    variable b1032 : boolean := false;
    variable b1031 : boolean := false;
    variable b1030 : boolean := false;
    variable b1029 : boolean := false;
    variable b1028 : boolean := false;
    variable b1027 : boolean := false;
    variable b1026 : boolean := false;
    variable r1025 : std_logic_vector(0 to 7) := (others => '0');
    variable r1024 : std_logic_vector(0 to 7) := (others => '0');
    variable r1023 : std_logic_vector(0 to 7) := (others => '0');
    variable r1022 : std_logic_vector(0 to 7) := (others => '0');
    variable r1021 : std_logic_vector(0 to 7) := (others => '0');
    variable r1020 : std_logic_vector(0 to 0) := (others => '0');
    variable r1019 : std_logic_vector(0 to 0) := (others => '0');
    variable r1018 : std_logic_vector(0 to 7) := (others => '0');
    variable r1017 : std_logic_vector(0 to 0) := (others => '0');
    variable r1016 : std_logic_vector(0 to 0) := (others => '0');
    variable r1015 : std_logic_vector(0 to 0) := (others => '0');
    variable r1014 : std_logic_vector(0 to 17) := (others => '0');
    variable r1013 : std_logic_vector(0 to 9) := (others => '0');
    variable b1012 : boolean := false;
    variable r1011 : std_logic_vector(0 to 7) := (others => '0');
  begin
    null;
    b1012 := true;
    r1013 := r1009(0 to 9);
    r1014 := r1009(10 to 27);
    r1015 := r1009(28 to 28);
    r1016 := r1009(29 to 29);
    r1017 := r1009(30 to 30);
    r1018 := r1009(31 to 38);
    r1019 := r1009(39 to 39);
    r1020 := r1009(40 to 40);
    r1021 := r1009(41 to 48);
    r1022 := r1009(49 to 56);
    r1023 := r1009(57 to 64);
    r1024 := r1009(65 to 72);
    r1025 := r1009(73 to 80);
    b1026 := true;
    b1027 := true;
    b1028 := true;
    b1029 := true;
    b1030 := true;
    b1031 := true;
    b1032 := true;
    b1033 := true;
    b1034 := true;
    b1035 := true;
    b1036 := true;
    b1037 := true;
    b1038 := true;
    b1039 := (b1026 AND (b1027 AND (b1028 AND (b1029 AND (b1030 AND (b1031 AND (b1032 AND (b1033 AND (b1034 AND (b1035 AND (b1036 AND (b1037 AND b1038))))))))))));
    if b1039 then
      null;
      r1011 := r1024;
    end if;
    return r1011;
  end rewire_r2_1008;
  function rewire_r1_969(r970 : std_logic_vector) return std_logic_vector
  is
    variable b1000 : boolean := false;
    variable b999 : boolean := false;
    variable b998 : boolean := false;
    variable b997 : boolean := false;
    variable b996 : boolean := false;
    variable b995 : boolean := false;
    variable b994 : boolean := false;
    variable b993 : boolean := false;
    variable b992 : boolean := false;
    variable b991 : boolean := false;
    variable b990 : boolean := false;
    variable b989 : boolean := false;
    variable b988 : boolean := false;
    variable b987 : boolean := false;
    variable r986 : std_logic_vector(0 to 7) := (others => '0');
    variable r985 : std_logic_vector(0 to 7) := (others => '0');
    variable r984 : std_logic_vector(0 to 7) := (others => '0');
    variable r983 : std_logic_vector(0 to 7) := (others => '0');
    variable r982 : std_logic_vector(0 to 7) := (others => '0');
    variable r981 : std_logic_vector(0 to 0) := (others => '0');
    variable r980 : std_logic_vector(0 to 0) := (others => '0');
    variable r979 : std_logic_vector(0 to 7) := (others => '0');
    variable r978 : std_logic_vector(0 to 0) := (others => '0');
    variable r977 : std_logic_vector(0 to 0) := (others => '0');
    variable r976 : std_logic_vector(0 to 0) := (others => '0');
    variable r975 : std_logic_vector(0 to 17) := (others => '0');
    variable r974 : std_logic_vector(0 to 9) := (others => '0');
    variable b973 : boolean := false;
    variable r972 : std_logic_vector(0 to 7) := (others => '0');
  begin
    null;
    b973 := true;
    r974 := r970(0 to 9);
    r975 := r970(10 to 27);
    r976 := r970(28 to 28);
    r977 := r970(29 to 29);
    r978 := r970(30 to 30);
    r979 := r970(31 to 38);
    r980 := r970(39 to 39);
    r981 := r970(40 to 40);
    r982 := r970(41 to 48);
    r983 := r970(49 to 56);
    r984 := r970(57 to 64);
    r985 := r970(65 to 72);
    r986 := r970(73 to 80);
    b987 := true;
    b988 := true;
    b989 := true;
    b990 := true;
    b991 := true;
    b992 := true;
    b993 := true;
    b994 := true;
    b995 := true;
    b996 := true;
    b997 := true;
    b998 := true;
    b999 := true;
    b1000 := (b987 AND (b988 AND (b989 AND (b990 AND (b991 AND (b992 AND (b993 AND (b994 AND (b995 AND (b996 AND (b997 AND (b998 AND b999))))))))))));
    if b1000 then
      null;
      r972 := r984;
    end if;
    return r972;
  end rewire_r1_969;
  function rewire_r0_930(r931 : std_logic_vector) return std_logic_vector
  is
    variable b961 : boolean := false;
    variable b960 : boolean := false;
    variable b959 : boolean := false;
    variable b958 : boolean := false;
    variable b957 : boolean := false;
    variable b956 : boolean := false;
    variable b955 : boolean := false;
    variable b954 : boolean := false;
    variable b953 : boolean := false;
    variable b952 : boolean := false;
    variable b951 : boolean := false;
    variable b950 : boolean := false;
    variable b949 : boolean := false;
    variable b948 : boolean := false;
    variable r947 : std_logic_vector(0 to 7) := (others => '0');
    variable r946 : std_logic_vector(0 to 7) := (others => '0');
    variable r945 : std_logic_vector(0 to 7) := (others => '0');
    variable r944 : std_logic_vector(0 to 7) := (others => '0');
    variable r943 : std_logic_vector(0 to 7) := (others => '0');
    variable r942 : std_logic_vector(0 to 0) := (others => '0');
    variable r941 : std_logic_vector(0 to 0) := (others => '0');
    variable r940 : std_logic_vector(0 to 7) := (others => '0');
    variable r939 : std_logic_vector(0 to 0) := (others => '0');
    variable r938 : std_logic_vector(0 to 0) := (others => '0');
    variable r937 : std_logic_vector(0 to 0) := (others => '0');
    variable r936 : std_logic_vector(0 to 17) := (others => '0');
    variable r935 : std_logic_vector(0 to 9) := (others => '0');
    variable b934 : boolean := false;
    variable r933 : std_logic_vector(0 to 7) := (others => '0');
  begin
    null;
    b934 := true;
    r935 := r931(0 to 9);
    r936 := r931(10 to 27);
    r937 := r931(28 to 28);
    r938 := r931(29 to 29);
    r939 := r931(30 to 30);
    r940 := r931(31 to 38);
    r941 := r931(39 to 39);
    r942 := r931(40 to 40);
    r943 := r931(41 to 48);
    r944 := r931(49 to 56);
    r945 := r931(57 to 64);
    r946 := r931(65 to 72);
    r947 := r931(73 to 80);
    b948 := true;
    b949 := true;
    b950 := true;
    b951 := true;
    b952 := true;
    b953 := true;
    b954 := true;
    b955 := true;
    b956 := true;
    b957 := true;
    b958 := true;
    b959 := true;
    b960 := true;
    b961 := (b948 AND (b949 AND (b950 AND (b951 AND (b952 AND (b953 AND (b954 AND (b955 AND (b956 AND (b957 AND (b958 AND (b959 AND b960))))))))))));
    if b961 then
      null;
      r933 := r944;
    end if;
    return r933;
  end rewire_r0_930;
  function rewire_mkReg_883(r884 : std_logic_vector ; r885 : std_logic_vector) return std_logic_vector
  is
    variable r920 : std_logic_vector(0 to 1) := (others => '0');
    variable b919 : boolean := false;
    variable b918 : boolean := false;
    variable b917 : boolean := false;
    variable r916 : std_logic_vector(0 to 0) := (others => '0');
    variable r915 : std_logic_vector(0 to 0) := (others => '0');
    variable b914 : boolean := false;
    variable r912 : std_logic_vector(0 to 1) := (others => '0');
    variable b911 : boolean := false;
    variable b910 : boolean := false;
    variable b909 : boolean := false;
    variable r908 : std_logic_vector(0 to 0) := (others => '0');
    variable r907 : std_logic_vector(0 to 0) := (others => '0');
    variable b906 : boolean := false;
    variable r904 : std_logic_vector(0 to 1) := (others => '0');
    variable b903 : boolean := false;
    variable b902 : boolean := false;
    variable b901 : boolean := false;
    variable r900 : std_logic_vector(0 to 0) := (others => '0');
    variable r899 : std_logic_vector(0 to 0) := (others => '0');
    variable b898 : boolean := false;
    variable r896 : std_logic_vector(0 to 1) := (others => '0');
    variable b895 : boolean := false;
    variable b894 : boolean := false;
    variable b893 : boolean := false;
    variable r892 : std_logic_vector(0 to 0) := (others => '0');
    variable r891 : std_logic_vector(0 to 0) := (others => '0');
    variable b890 : boolean := false;
    variable r889 : std_logic_vector(0 to 1) := (others => '0');
    variable r888 : std_logic_vector(0 to 1) := (others => '0');
    variable EMPTY : std_logic_vector(0 to -1) := (others => '0');
  begin
    null;
    null;
    r888 := (r884 & r885);
    b890 := true;
    r891 := r888(0 to 0);
    r892 := r888(1 to 1);
    b893 := ("0" = r891(0 to 0));
    b894 := ("0" = r892(0 to 0));
    b895 := (b893 AND b894);
    if b895 then
      r896 := "00";
      r889 := r896;
    end if;
    b898 := true;
    r899 := r888(0 to 0);
    r900 := r888(1 to 1);
    b901 := ("0" = r899(0 to 0));
    b902 := ("1" = r900(0 to 0));
    b903 := (b901 AND b902);
    if b903 then
      r904 := "01";
      r889 := r904;
    end if;
    b906 := true;
    r907 := r888(0 to 0);
    r908 := r888(1 to 1);
    b909 := ("1" = r907(0 to 0));
    b910 := ("0" = r908(0 to 0));
    b911 := (b909 AND b910);
    if b911 then
      r912 := "10";
      r889 := r912;
    end if;
    b914 := true;
    r915 := r888(0 to 0);
    r916 := r888(1 to 1);
    b917 := ("1" = r915(0 to 0));
    b918 := ("1" = r916(0 to 0));
    b919 := (b917 AND b918);
    if b919 then
      r920 := "11";
      r889 := r920;
    end if;
    return r889;
  end rewire_mkReg_883;
  function rewire_setWeOut_853(r854 : std_logic_vector ; r855 : std_logic_vector) return std_logic_vector
  is
    variable r869 : std_logic_vector(0 to 17) := (others => '0');
    variable EMPTY : std_logic_vector(0 to -1) := (others => '0');
    variable b867 : boolean := false;
    variable b866 : boolean := false;
    variable b865 : boolean := false;
    variable b864 : boolean := false;
    variable b863 : boolean := false;
    variable r862 : std_logic_vector(0 to 0) := (others => '0');
    variable r861 : std_logic_vector(0 to 0) := (others => '0');
    variable r860 : std_logic_vector(0 to 7) := (others => '0');
    variable r859 : std_logic_vector(0 to 7) := (others => '0');
    variable b858 : boolean := false;
    variable r857 : std_logic_vector(0 to 17) := (others => '0');
  begin
    null;
    b858 := true;
    r859 := r854(0 to 7);
    r860 := r854(8 to 15);
    r861 := r854(16 to 16);
    r862 := r854(17 to 17);
    b863 := true;
    b864 := true;
    b865 := true;
    b866 := true;
    b867 := (b863 AND (b864 AND (b865 AND b866)));
    if b867 then
      null;
      null;
      null;
      null;
      r869 := (r859 & r860 & r855 & r862);
      r857 := r869;
    end if;
    return r857;
  end rewire_setWeOut_853;
  function rewire_setAddrOut_782(r783 : std_logic_vector ; r784 : std_logic_vector) return std_logic_vector
  is
    variable r798 : std_logic_vector(0 to 17) := (others => '0');
    variable EMPTY : std_logic_vector(0 to -1) := (others => '0');
    variable b796 : boolean := false;
    variable b795 : boolean := false;
    variable b794 : boolean := false;
    variable b793 : boolean := false;
    variable b792 : boolean := false;
    variable r791 : std_logic_vector(0 to 0) := (others => '0');
    variable r790 : std_logic_vector(0 to 0) := (others => '0');
    variable r789 : std_logic_vector(0 to 7) := (others => '0');
    variable r788 : std_logic_vector(0 to 7) := (others => '0');
    variable b787 : boolean := false;
    variable r786 : std_logic_vector(0 to 17) := (others => '0');
  begin
    null;
    b787 := true;
    r788 := r783(0 to 7);
    r789 := r783(8 to 15);
    r790 := r783(16 to 16);
    r791 := r783(17 to 17);
    b792 := true;
    b793 := true;
    b794 := true;
    b795 := true;
    b796 := (b792 AND (b793 AND (b794 AND b795)));
    if b796 then
      null;
      null;
      null;
      null;
      r798 := (r784 & r789 & r790 & r791);
      r786 := r798;
    end if;
    return r786;
  end rewire_setAddrOut_782;
  function rewire_dataIn_717(r718 : std_logic_vector) return std_logic_vector
  is
    variable b728 : boolean := false;
    variable b727 : boolean := false;
    variable b726 : boolean := false;
    variable b725 : boolean := false;
    variable r724 : std_logic_vector(0 to 0) := (others => '0');
    variable r723 : std_logic_vector(0 to 0) := (others => '0');
    variable r722 : std_logic_vector(0 to 7) := (others => '0');
    variable b721 : boolean := false;
    variable r720 : std_logic_vector(0 to 7) := (others => '0');
  begin
    null;
    b721 := true;
    r722 := r718(0 to 7);
    r723 := r718(8 to 8);
    r724 := r718(9 to 9);
    b725 := true;
    b726 := true;
    b727 := true;
    b728 := (b725 AND (b726 AND b727));
    if b728 then
      null;
      r720 := r722;
    end if;
    return r720;
  end rewire_dataIn_717;
  function rewire_setCSave_657(r658 : std_logic_vector ; r659 : std_logic_vector) return std_logic_vector
  is
    variable r691 : std_logic_vector(0 to 80) := (others => '0');
    variable EMPTY : std_logic_vector(0 to -1) := (others => '0');
    variable b689 : boolean := false;
    variable b688 : boolean := false;
    variable b687 : boolean := false;
    variable b686 : boolean := false;
    variable b685 : boolean := false;
    variable b684 : boolean := false;
    variable b683 : boolean := false;
    variable b682 : boolean := false;
    variable b681 : boolean := false;
    variable b680 : boolean := false;
    variable b679 : boolean := false;
    variable b678 : boolean := false;
    variable b677 : boolean := false;
    variable b676 : boolean := false;
    variable r675 : std_logic_vector(0 to 7) := (others => '0');
    variable r674 : std_logic_vector(0 to 7) := (others => '0');
    variable r673 : std_logic_vector(0 to 7) := (others => '0');
    variable r672 : std_logic_vector(0 to 7) := (others => '0');
    variable r671 : std_logic_vector(0 to 7) := (others => '0');
    variable r670 : std_logic_vector(0 to 0) := (others => '0');
    variable r669 : std_logic_vector(0 to 0) := (others => '0');
    variable r668 : std_logic_vector(0 to 7) := (others => '0');
    variable r667 : std_logic_vector(0 to 0) := (others => '0');
    variable r666 : std_logic_vector(0 to 0) := (others => '0');
    variable r665 : std_logic_vector(0 to 0) := (others => '0');
    variable r664 : std_logic_vector(0 to 17) := (others => '0');
    variable r663 : std_logic_vector(0 to 9) := (others => '0');
    variable b662 : boolean := false;
    variable r661 : std_logic_vector(0 to 80) := (others => '0');
  begin
    null;
    b662 := true;
    r663 := r658(0 to 9);
    r664 := r658(10 to 27);
    r665 := r658(28 to 28);
    r666 := r658(29 to 29);
    r667 := r658(30 to 30);
    r668 := r658(31 to 38);
    r669 := r658(39 to 39);
    r670 := r658(40 to 40);
    r671 := r658(41 to 48);
    r672 := r658(49 to 56);
    r673 := r658(57 to 64);
    r674 := r658(65 to 72);
    r675 := r658(73 to 80);
    b676 := true;
    b677 := true;
    b678 := true;
    b679 := true;
    b680 := true;
    b681 := true;
    b682 := true;
    b683 := true;
    b684 := true;
    b685 := true;
    b686 := true;
    b687 := true;
    b688 := true;
    b689 := (b676 AND (b677 AND (b678 AND (b679 AND (b680 AND (b681 AND (b682 AND (b683 AND (b684 AND (b685 AND (b686 AND (b687 AND b688))))))))))));
    if b689 then
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      r691 := (r663 & r664 & r665 & r666 & r667 & r668 & r669 & r659 & r671 & r672 & r673 & r674 & r675);
      r661 := r691;
    end if;
    return r661;
  end rewire_setCSave_657;
  function rewire_setZSave_615(r616 : std_logic_vector ; r617 : std_logic_vector) return std_logic_vector
  is
    variable r649 : std_logic_vector(0 to 80) := (others => '0');
    variable EMPTY : std_logic_vector(0 to -1) := (others => '0');
    variable b647 : boolean := false;
    variable b646 : boolean := false;
    variable b645 : boolean := false;
    variable b644 : boolean := false;
    variable b643 : boolean := false;
    variable b642 : boolean := false;
    variable b641 : boolean := false;
    variable b640 : boolean := false;
    variable b639 : boolean := false;
    variable b638 : boolean := false;
    variable b637 : boolean := false;
    variable b636 : boolean := false;
    variable b635 : boolean := false;
    variable b634 : boolean := false;
    variable r633 : std_logic_vector(0 to 7) := (others => '0');
    variable r632 : std_logic_vector(0 to 7) := (others => '0');
    variable r631 : std_logic_vector(0 to 7) := (others => '0');
    variable r630 : std_logic_vector(0 to 7) := (others => '0');
    variable r629 : std_logic_vector(0 to 7) := (others => '0');
    variable r628 : std_logic_vector(0 to 0) := (others => '0');
    variable r627 : std_logic_vector(0 to 0) := (others => '0');
    variable r626 : std_logic_vector(0 to 7) := (others => '0');
    variable r625 : std_logic_vector(0 to 0) := (others => '0');
    variable r624 : std_logic_vector(0 to 0) := (others => '0');
    variable r623 : std_logic_vector(0 to 0) := (others => '0');
    variable r622 : std_logic_vector(0 to 17) := (others => '0');
    variable r621 : std_logic_vector(0 to 9) := (others => '0');
    variable b620 : boolean := false;
    variable r619 : std_logic_vector(0 to 80) := (others => '0');
  begin
    null;
    b620 := true;
    r621 := r616(0 to 9);
    r622 := r616(10 to 27);
    r623 := r616(28 to 28);
    r624 := r616(29 to 29);
    r625 := r616(30 to 30);
    r626 := r616(31 to 38);
    r627 := r616(39 to 39);
    r628 := r616(40 to 40);
    r629 := r616(41 to 48);
    r630 := r616(49 to 56);
    r631 := r616(57 to 64);
    r632 := r616(65 to 72);
    r633 := r616(73 to 80);
    b634 := true;
    b635 := true;
    b636 := true;
    b637 := true;
    b638 := true;
    b639 := true;
    b640 := true;
    b641 := true;
    b642 := true;
    b643 := true;
    b644 := true;
    b645 := true;
    b646 := true;
    b647 := (b634 AND (b635 AND (b636 AND (b637 AND (b638 AND (b639 AND (b640 AND (b641 AND (b642 AND (b643 AND (b644 AND (b645 AND b646))))))))))));
    if b647 then
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      r649 := (r621 & r622 & r623 & r624 & r625 & r626 & r617 & r628 & r629 & r630 & r631 & r632 & r633);
      r619 := r649;
    end if;
    return r619;
  end rewire_setZSave_615;
  function rewire_setPCSave_573(r574 : std_logic_vector ; r575 : std_logic_vector) return std_logic_vector
  is
    variable r607 : std_logic_vector(0 to 80) := (others => '0');
    variable EMPTY : std_logic_vector(0 to -1) := (others => '0');
    variable b605 : boolean := false;
    variable b604 : boolean := false;
    variable b603 : boolean := false;
    variable b602 : boolean := false;
    variable b601 : boolean := false;
    variable b600 : boolean := false;
    variable b599 : boolean := false;
    variable b598 : boolean := false;
    variable b597 : boolean := false;
    variable b596 : boolean := false;
    variable b595 : boolean := false;
    variable b594 : boolean := false;
    variable b593 : boolean := false;
    variable b592 : boolean := false;
    variable r591 : std_logic_vector(0 to 7) := (others => '0');
    variable r590 : std_logic_vector(0 to 7) := (others => '0');
    variable r589 : std_logic_vector(0 to 7) := (others => '0');
    variable r588 : std_logic_vector(0 to 7) := (others => '0');
    variable r587 : std_logic_vector(0 to 7) := (others => '0');
    variable r586 : std_logic_vector(0 to 0) := (others => '0');
    variable r585 : std_logic_vector(0 to 0) := (others => '0');
    variable r584 : std_logic_vector(0 to 7) := (others => '0');
    variable r583 : std_logic_vector(0 to 0) := (others => '0');
    variable r582 : std_logic_vector(0 to 0) := (others => '0');
    variable r581 : std_logic_vector(0 to 0) := (others => '0');
    variable r580 : std_logic_vector(0 to 17) := (others => '0');
    variable r579 : std_logic_vector(0 to 9) := (others => '0');
    variable b578 : boolean := false;
    variable r577 : std_logic_vector(0 to 80) := (others => '0');
  begin
    null;
    b578 := true;
    r579 := r574(0 to 9);
    r580 := r574(10 to 27);
    r581 := r574(28 to 28);
    r582 := r574(29 to 29);
    r583 := r574(30 to 30);
    r584 := r574(31 to 38);
    r585 := r574(39 to 39);
    r586 := r574(40 to 40);
    r587 := r574(41 to 48);
    r588 := r574(49 to 56);
    r589 := r574(57 to 64);
    r590 := r574(65 to 72);
    r591 := r574(73 to 80);
    b592 := true;
    b593 := true;
    b594 := true;
    b595 := true;
    b596 := true;
    b597 := true;
    b598 := true;
    b599 := true;
    b600 := true;
    b601 := true;
    b602 := true;
    b603 := true;
    b604 := true;
    b605 := (b592 AND (b593 AND (b594 AND (b595 AND (b596 AND (b597 AND (b598 AND (b599 AND (b600 AND (b601 AND (b602 AND (b603 AND b604))))))))))));
    if b605 then
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      r607 := (r579 & r580 & r581 & r582 & r583 & r584 & r585 & r586 & r575 & r588 & r589 & r590 & r591);
      r577 := r607;
    end if;
    return r577;
  end rewire_setPCSave_573;
  function rewire_cFlag_536(r537 : std_logic_vector) return std_logic_vector
  is
    variable b567 : boolean := false;
    variable b566 : boolean := false;
    variable b565 : boolean := false;
    variable b564 : boolean := false;
    variable b563 : boolean := false;
    variable b562 : boolean := false;
    variable b561 : boolean := false;
    variable b560 : boolean := false;
    variable b559 : boolean := false;
    variable b558 : boolean := false;
    variable b557 : boolean := false;
    variable b556 : boolean := false;
    variable b555 : boolean := false;
    variable b554 : boolean := false;
    variable r553 : std_logic_vector(0 to 7) := (others => '0');
    variable r552 : std_logic_vector(0 to 7) := (others => '0');
    variable r551 : std_logic_vector(0 to 7) := (others => '0');
    variable r550 : std_logic_vector(0 to 7) := (others => '0');
    variable r549 : std_logic_vector(0 to 7) := (others => '0');
    variable r548 : std_logic_vector(0 to 0) := (others => '0');
    variable r547 : std_logic_vector(0 to 0) := (others => '0');
    variable r546 : std_logic_vector(0 to 7) := (others => '0');
    variable r545 : std_logic_vector(0 to 0) := (others => '0');
    variable r544 : std_logic_vector(0 to 0) := (others => '0');
    variable r543 : std_logic_vector(0 to 0) := (others => '0');
    variable r542 : std_logic_vector(0 to 17) := (others => '0');
    variable r541 : std_logic_vector(0 to 9) := (others => '0');
    variable b540 : boolean := false;
    variable r539 : std_logic_vector(0 to 0) := (others => '0');
  begin
    null;
    b540 := true;
    r541 := r537(0 to 9);
    r542 := r537(10 to 27);
    r543 := r537(28 to 28);
    r544 := r537(29 to 29);
    r545 := r537(30 to 30);
    r546 := r537(31 to 38);
    r547 := r537(39 to 39);
    r548 := r537(40 to 40);
    r549 := r537(41 to 48);
    r550 := r537(49 to 56);
    r551 := r537(57 to 64);
    r552 := r537(65 to 72);
    r553 := r537(73 to 80);
    b554 := true;
    b555 := true;
    b556 := true;
    b557 := true;
    b558 := true;
    b559 := true;
    b560 := true;
    b561 := true;
    b562 := true;
    b563 := true;
    b564 := true;
    b565 := true;
    b566 := true;
    b567 := (b554 AND (b555 AND (b556 AND (b557 AND (b558 AND (b559 AND (b560 AND (b561 AND (b562 AND (b563 AND (b564 AND (b565 AND b566))))))))))));
    if b567 then
      null;
      r539 := r544;
    end if;
    return r539;
  end rewire_cFlag_536;
  function rewire_zFlag_499(r500 : std_logic_vector) return std_logic_vector
  is
    variable b530 : boolean := false;
    variable b529 : boolean := false;
    variable b528 : boolean := false;
    variable b527 : boolean := false;
    variable b526 : boolean := false;
    variable b525 : boolean := false;
    variable b524 : boolean := false;
    variable b523 : boolean := false;
    variable b522 : boolean := false;
    variable b521 : boolean := false;
    variable b520 : boolean := false;
    variable b519 : boolean := false;
    variable b518 : boolean := false;
    variable b517 : boolean := false;
    variable r516 : std_logic_vector(0 to 7) := (others => '0');
    variable r515 : std_logic_vector(0 to 7) := (others => '0');
    variable r514 : std_logic_vector(0 to 7) := (others => '0');
    variable r513 : std_logic_vector(0 to 7) := (others => '0');
    variable r512 : std_logic_vector(0 to 7) := (others => '0');
    variable r511 : std_logic_vector(0 to 0) := (others => '0');
    variable r510 : std_logic_vector(0 to 0) := (others => '0');
    variable r509 : std_logic_vector(0 to 7) := (others => '0');
    variable r508 : std_logic_vector(0 to 0) := (others => '0');
    variable r507 : std_logic_vector(0 to 0) := (others => '0');
    variable r506 : std_logic_vector(0 to 0) := (others => '0');
    variable r505 : std_logic_vector(0 to 17) := (others => '0');
    variable r504 : std_logic_vector(0 to 9) := (others => '0');
    variable b503 : boolean := false;
    variable r502 : std_logic_vector(0 to 0) := (others => '0');
  begin
    null;
    b503 := true;
    r504 := r500(0 to 9);
    r505 := r500(10 to 27);
    r506 := r500(28 to 28);
    r507 := r500(29 to 29);
    r508 := r500(30 to 30);
    r509 := r500(31 to 38);
    r510 := r500(39 to 39);
    r511 := r500(40 to 40);
    r512 := r500(41 to 48);
    r513 := r500(49 to 56);
    r514 := r500(57 to 64);
    r515 := r500(65 to 72);
    r516 := r500(73 to 80);
    b517 := true;
    b518 := true;
    b519 := true;
    b520 := true;
    b521 := true;
    b522 := true;
    b523 := true;
    b524 := true;
    b525 := true;
    b526 := true;
    b527 := true;
    b528 := true;
    b529 := true;
    b530 := (b517 AND (b518 AND (b519 AND (b520 AND (b521 AND (b522 AND (b523 AND (b524 AND (b525 AND (b526 AND (b527 AND (b528 AND b529))))))))))));
    if b530 then
      null;
      r502 := r506;
    end if;
    return r502;
  end rewire_zFlag_499;
  function rewire_pc_462(r463 : std_logic_vector) return std_logic_vector
  is
    variable b493 : boolean := false;
    variable b492 : boolean := false;
    variable b491 : boolean := false;
    variable b490 : boolean := false;
    variable b489 : boolean := false;
    variable b488 : boolean := false;
    variable b487 : boolean := false;
    variable b486 : boolean := false;
    variable b485 : boolean := false;
    variable b484 : boolean := false;
    variable b483 : boolean := false;
    variable b482 : boolean := false;
    variable b481 : boolean := false;
    variable b480 : boolean := false;
    variable r479 : std_logic_vector(0 to 7) := (others => '0');
    variable r478 : std_logic_vector(0 to 7) := (others => '0');
    variable r477 : std_logic_vector(0 to 7) := (others => '0');
    variable r476 : std_logic_vector(0 to 7) := (others => '0');
    variable r475 : std_logic_vector(0 to 7) := (others => '0');
    variable r474 : std_logic_vector(0 to 0) := (others => '0');
    variable r473 : std_logic_vector(0 to 0) := (others => '0');
    variable r472 : std_logic_vector(0 to 7) := (others => '0');
    variable r471 : std_logic_vector(0 to 0) := (others => '0');
    variable r470 : std_logic_vector(0 to 0) := (others => '0');
    variable r469 : std_logic_vector(0 to 0) := (others => '0');
    variable r468 : std_logic_vector(0 to 17) := (others => '0');
    variable r467 : std_logic_vector(0 to 9) := (others => '0');
    variable b466 : boolean := false;
    variable r465 : std_logic_vector(0 to 7) := (others => '0');
  begin
    null;
    b466 := true;
    r467 := r463(0 to 9);
    r468 := r463(10 to 27);
    r469 := r463(28 to 28);
    r470 := r463(29 to 29);
    r471 := r463(30 to 30);
    r472 := r463(31 to 38);
    r473 := r463(39 to 39);
    r474 := r463(40 to 40);
    r475 := r463(41 to 48);
    r476 := r463(49 to 56);
    r477 := r463(57 to 64);
    r478 := r463(65 to 72);
    r479 := r463(73 to 80);
    b480 := true;
    b481 := true;
    b482 := true;
    b483 := true;
    b484 := true;
    b485 := true;
    b486 := true;
    b487 := true;
    b488 := true;
    b489 := true;
    b490 := true;
    b491 := true;
    b492 := true;
    b493 := (b480 AND (b481 AND (b482 AND (b483 AND (b484 AND (b485 AND (b486 AND (b487 AND (b488 AND (b489 AND (b490 AND (b491 AND b492))))))))))));
    if b493 then
      null;
      r465 := r472;
    end if;
    return r465;
  end rewire_pc_462;
  function rewire_setIEFlag_419(r420 : std_logic_vector ; r421 : std_logic_vector) return std_logic_vector
  is
    variable r453 : std_logic_vector(0 to 80) := (others => '0');
    variable EMPTY : std_logic_vector(0 to -1) := (others => '0');
    variable b451 : boolean := false;
    variable b450 : boolean := false;
    variable b449 : boolean := false;
    variable b448 : boolean := false;
    variable b447 : boolean := false;
    variable b446 : boolean := false;
    variable b445 : boolean := false;
    variable b444 : boolean := false;
    variable b443 : boolean := false;
    variable b442 : boolean := false;
    variable b441 : boolean := false;
    variable b440 : boolean := false;
    variable b439 : boolean := false;
    variable b438 : boolean := false;
    variable r437 : std_logic_vector(0 to 7) := (others => '0');
    variable r436 : std_logic_vector(0 to 7) := (others => '0');
    variable r435 : std_logic_vector(0 to 7) := (others => '0');
    variable r434 : std_logic_vector(0 to 7) := (others => '0');
    variable r433 : std_logic_vector(0 to 7) := (others => '0');
    variable r432 : std_logic_vector(0 to 0) := (others => '0');
    variable r431 : std_logic_vector(0 to 0) := (others => '0');
    variable r430 : std_logic_vector(0 to 7) := (others => '0');
    variable r429 : std_logic_vector(0 to 0) := (others => '0');
    variable r428 : std_logic_vector(0 to 0) := (others => '0');
    variable r427 : std_logic_vector(0 to 0) := (others => '0');
    variable r426 : std_logic_vector(0 to 17) := (others => '0');
    variable r425 : std_logic_vector(0 to 9) := (others => '0');
    variable b424 : boolean := false;
    variable r423 : std_logic_vector(0 to 80) := (others => '0');
  begin
    null;
    b424 := true;
    r425 := r420(0 to 9);
    r426 := r420(10 to 27);
    r427 := r420(28 to 28);
    r428 := r420(29 to 29);
    r429 := r420(30 to 30);
    r430 := r420(31 to 38);
    r431 := r420(39 to 39);
    r432 := r420(40 to 40);
    r433 := r420(41 to 48);
    r434 := r420(49 to 56);
    r435 := r420(57 to 64);
    r436 := r420(65 to 72);
    r437 := r420(73 to 80);
    b438 := true;
    b439 := true;
    b440 := true;
    b441 := true;
    b442 := true;
    b443 := true;
    b444 := true;
    b445 := true;
    b446 := true;
    b447 := true;
    b448 := true;
    b449 := true;
    b450 := true;
    b451 := (b438 AND (b439 AND (b440 AND (b441 AND (b442 AND (b443 AND (b444 AND (b445 AND (b446 AND (b447 AND (b448 AND (b449 AND b450))))))))))));
    if b451 then
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      r453 := (r425 & r426 & r427 & r428 & r421 & r430 & r431 & r432 & r433 & r434 & r435 & r436 & r437);
      r423 := r453;
    end if;
    return r423;
  end rewire_setIEFlag_419;
  function rewire_intIn_387(r388 : std_logic_vector) return std_logic_vector
  is
    variable b398 : boolean := false;
    variable b397 : boolean := false;
    variable b396 : boolean := false;
    variable b395 : boolean := false;
    variable r394 : std_logic_vector(0 to 0) := (others => '0');
    variable r393 : std_logic_vector(0 to 0) := (others => '0');
    variable r392 : std_logic_vector(0 to 7) := (others => '0');
    variable b391 : boolean := false;
    variable r390 : std_logic_vector(0 to 0) := (others => '0');
  begin
    null;
    b391 := true;
    r392 := r388(0 to 7);
    r393 := r388(8 to 8);
    r394 := r388(9 to 9);
    b395 := true;
    b396 := true;
    b397 := true;
    b398 := (b395 AND (b396 AND b397));
    if b398 then
      null;
      r390 := r394;
    end if;
    return r390;
  end rewire_intIn_387;
  function rewire_rstIn_264(r265 : std_logic_vector) return std_logic_vector
  is
    variable b275 : boolean := false;
    variable b274 : boolean := false;
    variable b273 : boolean := false;
    variable b272 : boolean := false;
    variable r271 : std_logic_vector(0 to 0) := (others => '0');
    variable r270 : std_logic_vector(0 to 0) := (others => '0');
    variable r269 : std_logic_vector(0 to 7) := (others => '0');
    variable b268 : boolean := false;
    variable r267 : std_logic_vector(0 to 0) := (others => '0');
  begin
    null;
    b268 := true;
    r269 := r265(0 to 7);
    r270 := r265(8 to 8);
    r271 := r265(9 to 9);
    b272 := true;
    b273 := true;
    b274 := true;
    b275 := (b272 AND (b273 AND b274));
    if b275 then
      null;
      r267 := r270;
    end if;
    return r267;
  end rewire_rstIn_264;
  function rewire_inputs_229(r230 : std_logic_vector) return std_logic_vector
  is
    variable b260 : boolean := false;
    variable b259 : boolean := false;
    variable b258 : boolean := false;
    variable b257 : boolean := false;
    variable b256 : boolean := false;
    variable b255 : boolean := false;
    variable b254 : boolean := false;
    variable b253 : boolean := false;
    variable b252 : boolean := false;
    variable b251 : boolean := false;
    variable b250 : boolean := false;
    variable b249 : boolean := false;
    variable b248 : boolean := false;
    variable b247 : boolean := false;
    variable r246 : std_logic_vector(0 to 7) := (others => '0');
    variable r245 : std_logic_vector(0 to 7) := (others => '0');
    variable r244 : std_logic_vector(0 to 7) := (others => '0');
    variable r243 : std_logic_vector(0 to 7) := (others => '0');
    variable r242 : std_logic_vector(0 to 7) := (others => '0');
    variable r241 : std_logic_vector(0 to 0) := (others => '0');
    variable r240 : std_logic_vector(0 to 0) := (others => '0');
    variable r239 : std_logic_vector(0 to 7) := (others => '0');
    variable r238 : std_logic_vector(0 to 0) := (others => '0');
    variable r237 : std_logic_vector(0 to 0) := (others => '0');
    variable r236 : std_logic_vector(0 to 0) := (others => '0');
    variable r235 : std_logic_vector(0 to 17) := (others => '0');
    variable r234 : std_logic_vector(0 to 9) := (others => '0');
    variable b233 : boolean := false;
    variable r232 : std_logic_vector(0 to 9) := (others => '0');
  begin
    null;
    b233 := true;
    r234 := r230(0 to 9);
    r235 := r230(10 to 27);
    r236 := r230(28 to 28);
    r237 := r230(29 to 29);
    r238 := r230(30 to 30);
    r239 := r230(31 to 38);
    r240 := r230(39 to 39);
    r241 := r230(40 to 40);
    r242 := r230(41 to 48);
    r243 := r230(49 to 56);
    r244 := r230(57 to 64);
    r245 := r230(65 to 72);
    r246 := r230(73 to 80);
    b247 := true;
    b248 := true;
    b249 := true;
    b250 := true;
    b251 := true;
    b252 := true;
    b253 := true;
    b254 := true;
    b255 := true;
    b256 := true;
    b257 := true;
    b258 := true;
    b259 := true;
    b260 := (b247 AND (b248 AND (b249 AND (b250 AND (b251 AND (b252 AND (b253 AND (b254 AND (b255 AND (b256 AND (b257 AND (b258 AND b259))))))))))));
    if b260 then
      null;
      r232 := r234;
    end if;
    return r232;
  end rewire_inputs_229;
  function rewire_setInputs_185(r186 : std_logic_vector ; r187 : std_logic_vector) return std_logic_vector
  is
    variable r219 : std_logic_vector(0 to 80) := (others => '0');
    variable EMPTY : std_logic_vector(0 to -1) := (others => '0');
    variable b217 : boolean := false;
    variable b216 : boolean := false;
    variable b215 : boolean := false;
    variable b214 : boolean := false;
    variable b213 : boolean := false;
    variable b212 : boolean := false;
    variable b211 : boolean := false;
    variable b210 : boolean := false;
    variable b209 : boolean := false;
    variable b208 : boolean := false;
    variable b207 : boolean := false;
    variable b206 : boolean := false;
    variable b205 : boolean := false;
    variable b204 : boolean := false;
    variable r203 : std_logic_vector(0 to 7) := (others => '0');
    variable r202 : std_logic_vector(0 to 7) := (others => '0');
    variable r201 : std_logic_vector(0 to 7) := (others => '0');
    variable r200 : std_logic_vector(0 to 7) := (others => '0');
    variable r199 : std_logic_vector(0 to 7) := (others => '0');
    variable r198 : std_logic_vector(0 to 0) := (others => '0');
    variable r197 : std_logic_vector(0 to 0) := (others => '0');
    variable r196 : std_logic_vector(0 to 7) := (others => '0');
    variable r195 : std_logic_vector(0 to 0) := (others => '0');
    variable r194 : std_logic_vector(0 to 0) := (others => '0');
    variable r193 : std_logic_vector(0 to 0) := (others => '0');
    variable r192 : std_logic_vector(0 to 17) := (others => '0');
    variable r191 : std_logic_vector(0 to 9) := (others => '0');
    variable b190 : boolean := false;
    variable r189 : std_logic_vector(0 to 80) := (others => '0');
  begin
    null;
    b190 := true;
    r191 := r186(0 to 9);
    r192 := r186(10 to 27);
    r193 := r186(28 to 28);
    r194 := r186(29 to 29);
    r195 := r186(30 to 30);
    r196 := r186(31 to 38);
    r197 := r186(39 to 39);
    r198 := r186(40 to 40);
    r199 := r186(41 to 48);
    r200 := r186(49 to 56);
    r201 := r186(57 to 64);
    r202 := r186(65 to 72);
    r203 := r186(73 to 80);
    b204 := true;
    b205 := true;
    b206 := true;
    b207 := true;
    b208 := true;
    b209 := true;
    b210 := true;
    b211 := true;
    b212 := true;
    b213 := true;
    b214 := true;
    b215 := true;
    b216 := true;
    b217 := (b204 AND (b205 AND (b206 AND (b207 AND (b208 AND (b209 AND (b210 AND (b211 AND (b212 AND (b213 AND (b214 AND (b215 AND b216))))))))))));
    if b217 then
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      r219 := (r187 & r192 & r193 & r194 & r195 & r196 & r197 & r198 & r199 & r200 & r201 & r202 & r203);
      r189 := r219;
    end if;
    return r189;
  end rewire_setInputs_185;
  function rewire_outputs_144(r145 : std_logic_vector) return std_logic_vector
  is
    variable b175 : boolean := false;
    variable b174 : boolean := false;
    variable b173 : boolean := false;
    variable b172 : boolean := false;
    variable b171 : boolean := false;
    variable b170 : boolean := false;
    variable b169 : boolean := false;
    variable b168 : boolean := false;
    variable b167 : boolean := false;
    variable b166 : boolean := false;
    variable b165 : boolean := false;
    variable b164 : boolean := false;
    variable b163 : boolean := false;
    variable b162 : boolean := false;
    variable r161 : std_logic_vector(0 to 7) := (others => '0');
    variable r160 : std_logic_vector(0 to 7) := (others => '0');
    variable r159 : std_logic_vector(0 to 7) := (others => '0');
    variable r158 : std_logic_vector(0 to 7) := (others => '0');
    variable r157 : std_logic_vector(0 to 7) := (others => '0');
    variable r156 : std_logic_vector(0 to 0) := (others => '0');
    variable r155 : std_logic_vector(0 to 0) := (others => '0');
    variable r154 : std_logic_vector(0 to 7) := (others => '0');
    variable r153 : std_logic_vector(0 to 0) := (others => '0');
    variable r152 : std_logic_vector(0 to 0) := (others => '0');
    variable r151 : std_logic_vector(0 to 0) := (others => '0');
    variable r150 : std_logic_vector(0 to 17) := (others => '0');
    variable r149 : std_logic_vector(0 to 9) := (others => '0');
    variable b148 : boolean := false;
    variable r147 : std_logic_vector(0 to 17) := (others => '0');
  begin
    null;
    b148 := true;
    r149 := r145(0 to 9);
    r150 := r145(10 to 27);
    r151 := r145(28 to 28);
    r152 := r145(29 to 29);
    r153 := r145(30 to 30);
    r154 := r145(31 to 38);
    r155 := r145(39 to 39);
    r156 := r145(40 to 40);
    r157 := r145(41 to 48);
    r158 := r145(49 to 56);
    r159 := r145(57 to 64);
    r160 := r145(65 to 72);
    r161 := r145(73 to 80);
    b162 := true;
    b163 := true;
    b164 := true;
    b165 := true;
    b166 := true;
    b167 := true;
    b168 := true;
    b169 := true;
    b170 := true;
    b171 := true;
    b172 := true;
    b173 := true;
    b174 := true;
    b175 := (b162 AND (b163 AND (b164 AND (b165 AND (b166 AND (b167 AND (b168 AND (b169 AND (b170 AND (b171 AND (b172 AND (b173 AND b174))))))))))));
    if b175 then
      null;
      r147 := r150;
    end if;
    return r147;
  end rewire_outputs_144;
  function rewire_initOutputs_127 return std_logic_vector
  is
    variable r136 : std_logic_vector(0 to 17) := (others => '0');
    variable r134 : std_logic_vector(0 to 0) := (others => '0');
    variable r132 : std_logic_vector(0 to 0) := (others => '0');
    variable r131 : std_logic_vector(0 to 7) := (others => '0');
    variable r130 : std_logic_vector(0 to 7) := (others => '0');
    variable EMPTY : std_logic_vector(0 to -1) := (others => '0');
  begin
    r130 := zeroW8;
    r131 := zeroW8;
    r132 := "0";
    r134 := "0";
    r136 := (r130 & r131 & r132 & r134);
    return r136;
  end rewire_initOutputs_127;
  function rewire_setOutputs_91(r92 : std_logic_vector ; r93 : std_logic_vector) return std_logic_vector
  is
    variable r125 : std_logic_vector(0 to 80) := (others => '0');
    variable EMPTY : std_logic_vector(0 to -1) := (others => '0');
    variable b123 : boolean := false;
    variable b122 : boolean := false;
    variable b121 : boolean := false;
    variable b120 : boolean := false;
    variable b119 : boolean := false;
    variable b118 : boolean := false;
    variable b117 : boolean := false;
    variable b116 : boolean := false;
    variable b115 : boolean := false;
    variable b114 : boolean := false;
    variable b113 : boolean := false;
    variable b112 : boolean := false;
    variable b111 : boolean := false;
    variable b110 : boolean := false;
    variable r109 : std_logic_vector(0 to 7) := (others => '0');
    variable r108 : std_logic_vector(0 to 7) := (others => '0');
    variable r107 : std_logic_vector(0 to 7) := (others => '0');
    variable r106 : std_logic_vector(0 to 7) := (others => '0');
    variable r105 : std_logic_vector(0 to 7) := (others => '0');
    variable r104 : std_logic_vector(0 to 0) := (others => '0');
    variable r103 : std_logic_vector(0 to 0) := (others => '0');
    variable r102 : std_logic_vector(0 to 7) := (others => '0');
    variable r101 : std_logic_vector(0 to 0) := (others => '0');
    variable r100 : std_logic_vector(0 to 0) := (others => '0');
    variable r99 : std_logic_vector(0 to 0) := (others => '0');
    variable r98 : std_logic_vector(0 to 17) := (others => '0');
    variable r97 : std_logic_vector(0 to 9) := (others => '0');
    variable b96 : boolean := false;
    variable r95 : std_logic_vector(0 to 80) := (others => '0');
  begin
    null;
    b96 := true;
    r97 := r92(0 to 9);
    r98 := r92(10 to 27);
    r99 := r92(28 to 28);
    r100 := r92(29 to 29);
    r101 := r92(30 to 30);
    r102 := r92(31 to 38);
    r103 := r92(39 to 39);
    r104 := r92(40 to 40);
    r105 := r92(41 to 48);
    r106 := r92(49 to 56);
    r107 := r92(57 to 64);
    r108 := r92(65 to 72);
    r109 := r92(73 to 80);
    b110 := true;
    b111 := true;
    b112 := true;
    b113 := true;
    b114 := true;
    b115 := true;
    b116 := true;
    b117 := true;
    b118 := true;
    b119 := true;
    b120 := true;
    b121 := true;
    b122 := true;
    b123 := (b110 AND (b111 AND (b112 AND (b113 AND (b114 AND (b115 AND (b116 AND (b117 AND (b118 AND (b119 AND (b120 AND (b121 AND b122))))))))))));
    if b123 then
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      r125 := (r97 & r93 & r99 & r100 & r101 & r102 & r103 & r104 & r105 & r106 & r107 & r108 & r109);
      r95 := r125;
    end if;
    return r95;
  end rewire_setOutputs_91;
  function rewire_setZFlag_48(r49 : std_logic_vector ; r50 : std_logic_vector) return std_logic_vector
  is
    variable r82 : std_logic_vector(0 to 80) := (others => '0');
    variable EMPTY : std_logic_vector(0 to -1) := (others => '0');
    variable b80 : boolean := false;
    variable b79 : boolean := false;
    variable b78 : boolean := false;
    variable b77 : boolean := false;
    variable b76 : boolean := false;
    variable b75 : boolean := false;
    variable b74 : boolean := false;
    variable b73 : boolean := false;
    variable b72 : boolean := false;
    variable b71 : boolean := false;
    variable b70 : boolean := false;
    variable b69 : boolean := false;
    variable b68 : boolean := false;
    variable b67 : boolean := false;
    variable r66 : std_logic_vector(0 to 7) := (others => '0');
    variable r65 : std_logic_vector(0 to 7) := (others => '0');
    variable r64 : std_logic_vector(0 to 7) := (others => '0');
    variable r63 : std_logic_vector(0 to 7) := (others => '0');
    variable r62 : std_logic_vector(0 to 7) := (others => '0');
    variable r61 : std_logic_vector(0 to 0) := (others => '0');
    variable r60 : std_logic_vector(0 to 0) := (others => '0');
    variable r59 : std_logic_vector(0 to 7) := (others => '0');
    variable r58 : std_logic_vector(0 to 0) := (others => '0');
    variable r57 : std_logic_vector(0 to 0) := (others => '0');
    variable r56 : std_logic_vector(0 to 0) := (others => '0');
    variable r55 : std_logic_vector(0 to 17) := (others => '0');
    variable r54 : std_logic_vector(0 to 9) := (others => '0');
    variable b53 : boolean := false;
    variable r52 : std_logic_vector(0 to 80) := (others => '0');
  begin
    null;
    b53 := true;
    r54 := r49(0 to 9);
    r55 := r49(10 to 27);
    r56 := r49(28 to 28);
    r57 := r49(29 to 29);
    r58 := r49(30 to 30);
    r59 := r49(31 to 38);
    r60 := r49(39 to 39);
    r61 := r49(40 to 40);
    r62 := r49(41 to 48);
    r63 := r49(49 to 56);
    r64 := r49(57 to 64);
    r65 := r49(65 to 72);
    r66 := r49(73 to 80);
    b67 := true;
    b68 := true;
    b69 := true;
    b70 := true;
    b71 := true;
    b72 := true;
    b73 := true;
    b74 := true;
    b75 := true;
    b76 := true;
    b77 := true;
    b78 := true;
    b79 := true;
    b80 := (b67 AND (b68 AND (b69 AND (b70 AND (b71 AND (b72 AND (b73 AND (b74 AND (b75 AND (b76 AND (b77 AND (b78 AND b79))))))))))));
    if b80 then
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      r82 := (r54 & r55 & r50 & r57 & r58 & r59 & r60 & r61 & r62 & r63 & r64 & r65 & r66);
      r52 := r82;
    end if;
    return r52;
  end rewire_setZFlag_48;
  function rewire_setCFlag_5(r6 : std_logic_vector ; r7 : std_logic_vector) return std_logic_vector
  is
    variable r39 : std_logic_vector(0 to 80) := (others => '0');
    variable EMPTY : std_logic_vector(0 to -1) := (others => '0');
    variable b37 : boolean := false;
    variable b36 : boolean := false;
    variable b35 : boolean := false;
    variable b34 : boolean := false;
    variable b33 : boolean := false;
    variable b32 : boolean := false;
    variable b31 : boolean := false;
    variable b30 : boolean := false;
    variable b29 : boolean := false;
    variable b28 : boolean := false;
    variable b27 : boolean := false;
    variable b26 : boolean := false;
    variable b25 : boolean := false;
    variable b24 : boolean := false;
    variable r23 : std_logic_vector(0 to 7) := (others => '0');
    variable r22 : std_logic_vector(0 to 7) := (others => '0');
    variable r21 : std_logic_vector(0 to 7) := (others => '0');
    variable r20 : std_logic_vector(0 to 7) := (others => '0');
    variable r19 : std_logic_vector(0 to 7) := (others => '0');
    variable r18 : std_logic_vector(0 to 0) := (others => '0');
    variable r17 : std_logic_vector(0 to 0) := (others => '0');
    variable r16 : std_logic_vector(0 to 7) := (others => '0');
    variable r15 : std_logic_vector(0 to 0) := (others => '0');
    variable r14 : std_logic_vector(0 to 0) := (others => '0');
    variable r13 : std_logic_vector(0 to 0) := (others => '0');
    variable r12 : std_logic_vector(0 to 17) := (others => '0');
    variable r11 : std_logic_vector(0 to 9) := (others => '0');
    variable b10 : boolean := false;
    variable r9 : std_logic_vector(0 to 80) := (others => '0');
  begin
    null;
    b10 := true;
    r11 := r6(0 to 9);
    r12 := r6(10 to 27);
    r13 := r6(28 to 28);
    r14 := r6(29 to 29);
    r15 := r6(30 to 30);
    r16 := r6(31 to 38);
    r17 := r6(39 to 39);
    r18 := r6(40 to 40);
    r19 := r6(41 to 48);
    r20 := r6(49 to 56);
    r21 := r6(57 to 64);
    r22 := r6(65 to 72);
    r23 := r6(73 to 80);
    b24 := true;
    b25 := true;
    b26 := true;
    b27 := true;
    b28 := true;
    b29 := true;
    b30 := true;
    b31 := true;
    b32 := true;
    b33 := true;
    b34 := true;
    b35 := true;
    b36 := true;
    b37 := (b24 AND (b25 AND (b26 AND (b27 AND (b28 AND (b29 AND (b30 AND (b31 AND (b32 AND (b33 AND (b34 AND (b35 AND b36))))))))))));
    if b37 then
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      r39 := (r11 & r12 & r13 & r7 & r15 & r16 & r17 & r18 & r19 & r20 & r21 & r22 & r23);
      r9 := r39;
    end if;
    return r9;
  end rewire_setCFlag_5;

begin
  process (clk)
    variable goto_L5438 : boolean := false;
    variable goto_L5427 : boolean := false;
    variable goto_L5383 : boolean := false;
    variable goto_L5128 : boolean := false;
    variable goto_L5026 : boolean := false;
    variable goto_L4932 : boolean := false;
    variable goto_L4885 : boolean := false;
    variable goto_L4703 : boolean := false;
    variable goto_L4521 : boolean := false;
    variable goto_L4422 : boolean := false;
    variable goto_L4285 : boolean := false;
    variable goto_L4091 : boolean := false;
    variable goto_L4004 : boolean := false;
    variable goto_L3943 : boolean := false;
    variable goto_L3848 : boolean := false;
    variable goto_L3737 : boolean := false;
    variable goto_L3628 : boolean := false;
    variable goto_L3517 : boolean := false;
    variable goto_L3408 : boolean := false;
    variable goto_L3234 : boolean := false;
    variable goto_L3048 : boolean := false;
    variable goto_L2862 : boolean := false;
    variable goto_L2676 : boolean := false;
    variable goto_L2547 : boolean := false;
    variable goto_L2339 : boolean := false;
    variable goto_L2135 : boolean := false;
    variable goto_L1927 : boolean := false;
    variable goto_L1723 : boolean := false;
    variable goto_L1506 : boolean := false;
    variable goto_L1537 : boolean := false;
    variable goto_L1546 : boolean := false;
    variable goto_L1555 : boolean := false;
    variable goto_L1549 : boolean := false;
    variable goto_L1540 : boolean := false;
    variable goto_L1531 : boolean := false;
    variable goto_L1528 : boolean := false;
    variable goto_L1189 : boolean := false;
    variable goto_L1391 : boolean := false;
    variable goto_L1202 : boolean := false;
    variable goto_L1259 : boolean := false;
    variable goto_L1303 : boolean := false;
    variable goto_L1347 : boolean := false;
    variable goto_L1341 : boolean := false;
    variable goto_L1297 : boolean := false;
    variable goto_L1253 : boolean := false;
    variable goto_L1215 : boolean := false;
    variable goto_L1198 : boolean := false;
    variable goto_L814 : boolean := false;
    variable goto_L1115 : boolean := false;
    variable goto_L882 : boolean := false;
    variable goto_L966 : boolean := false;
    variable goto_L1005 : boolean := false;
    variable goto_L1044 : boolean := false;
    variable goto_L1040 : boolean := false;
    variable goto_L1001 : boolean := false;
    variable goto_L962 : boolean := false;
    variable goto_L927 : boolean := false;
    variable goto_L878 : boolean := false;
    variable goto_L732 : boolean := false;
    variable goto_L705 : boolean := false;
    variable goto_L404 : boolean := false;
    variable goto_L314 : boolean := false;
    variable goto_L279 : boolean := false;
    variable goto_L182 : boolean := false;
    variable goto_L225 : boolean := false;
    variable goto_L323 : boolean := false;
    variable goto_L714 : boolean := false;
    variable goto_L1396 : boolean := false;
    variable goto_L1564 : boolean := false;
    variable goto_L1732 : boolean := false;
    variable goto_L1936 : boolean := false;
    variable goto_L2144 : boolean := false;
    variable goto_L2348 : boolean := false;
    variable goto_L2556 : boolean := false;
    variable goto_L2685 : boolean := false;
    variable goto_L2871 : boolean := false;
    variable goto_L3057 : boolean := false;
    variable goto_L3243 : boolean := false;
    variable goto_L3417 : boolean := false;
    variable goto_L3526 : boolean := false;
    variable goto_L3637 : boolean := false;
    variable goto_L3746 : boolean := false;
    variable goto_L3857 : boolean := false;
    variable goto_L3952 : boolean := false;
    variable goto_L4013 : boolean := false;
    variable goto_L4100 : boolean := false;
    variable goto_L4294 : boolean := false;
    variable goto_L4431 : boolean := false;
    variable goto_L4530 : boolean := false;
    variable goto_L4712 : boolean := false;
    variable goto_L4894 : boolean := false;
    variable goto_L5138 : boolean := false;
    variable goto_L5392 : boolean := false;
    variable goto_L5176 : boolean := false;
    variable goto_L5189 : boolean := false;
    variable goto_L5196 : boolean := false;
    variable goto_L5203 : boolean := false;
    variable goto_L5199 : boolean := false;
    variable goto_L5192 : boolean := false;
    variable goto_L5185 : boolean := false;
    variable goto_L5182 : boolean := false;
    variable goto_L5234 : boolean := false;
    variable goto_L5253 : boolean := false;
    variable goto_L5273 : boolean := false;
    variable goto_L5266 : boolean := false;
    variable goto_L5247 : boolean := false;
    variable goto_L5227 : boolean := false;
    variable goto_L5287 : boolean := false;
    variable goto_L5331 : boolean := false;
    variable goto_L5340 : boolean := false;
    variable goto_L5349 : boolean := false;
    variable goto_L5343 : boolean := false;
    variable goto_L5334 : boolean := false;
    variable goto_L5325 : boolean := false;
    variable goto_L5322 : boolean := false;
    variable goto_L4931 : boolean := false;
    variable goto_L5035 : boolean := false;
    variable goto_L5051 : boolean := false;
    variable goto_L5058 : boolean := false;
    variable goto_L5065 : boolean := false;
    variable goto_L5061 : boolean := false;
    variable goto_L5054 : boolean := false;
    variable goto_L5047 : boolean := false;
    variable goto_L5044 : boolean := false;
    variable goto_L5088 : boolean := false;
    variable goto_L5099 : boolean := false;
    variable goto_L5110 : boolean := false;
    variable goto_L5102 : boolean := false;
    variable goto_L5091 : boolean := false;
    variable goto_L5080 : boolean := false;
    variable goto_L5077 : boolean := false;
    variable goto_L4936 : boolean := false;
    variable goto_L4949 : boolean := false;
    variable goto_L4956 : boolean := false;
    variable goto_L4963 : boolean := false;
    variable goto_L4959 : boolean := false;
    variable goto_L4952 : boolean := false;
    variable goto_L4945 : boolean := false;
    variable goto_L4942 : boolean := false;
    variable goto_L4986 : boolean := false;
    variable goto_L4997 : boolean := false;
    variable goto_L5008 : boolean := false;
    variable goto_L5000 : boolean := false;
    variable goto_L4989 : boolean := false;
    variable goto_L4978 : boolean := false;
    variable goto_L4975 : boolean := false;
    variable goto_L4750 : boolean := false;
    variable goto_L4763 : boolean := false;
    variable goto_L4770 : boolean := false;
    variable goto_L4777 : boolean := false;
    variable goto_L4773 : boolean := false;
    variable goto_L4766 : boolean := false;
    variable goto_L4759 : boolean := false;
    variable goto_L4756 : boolean := false;
    variable goto_L4833 : boolean := false;
    variable goto_L4842 : boolean := false;
    variable goto_L4851 : boolean := false;
    variable goto_L4845 : boolean := false;
    variable goto_L4836 : boolean := false;
    variable goto_L4827 : boolean := false;
    variable goto_L4824 : boolean := false;
    variable goto_L4568 : boolean := false;
    variable goto_L4581 : boolean := false;
    variable goto_L4588 : boolean := false;
    variable goto_L4595 : boolean := false;
    variable goto_L4591 : boolean := false;
    variable goto_L4584 : boolean := false;
    variable goto_L4577 : boolean := false;
    variable goto_L4574 : boolean := false;
    variable goto_L4651 : boolean := false;
    variable goto_L4660 : boolean := false;
    variable goto_L4669 : boolean := false;
    variable goto_L4663 : boolean := false;
    variable goto_L4654 : boolean := false;
    variable goto_L4645 : boolean := false;
    variable goto_L4642 : boolean := false;
    variable goto_L4469 : boolean := false;
    variable goto_L4484 : boolean := false;
    variable goto_L4494 : boolean := false;
    variable goto_L4504 : boolean := false;
    variable goto_L4497 : boolean := false;
    variable goto_L4487 : boolean := false;
    variable goto_L4477 : boolean := false;
    variable goto_L4474 : boolean := false;
    variable goto_L4332 : boolean := false;
    variable goto_L4345 : boolean := false;
    variable goto_L4352 : boolean := false;
    variable goto_L4359 : boolean := false;
    variable goto_L4355 : boolean := false;
    variable goto_L4348 : boolean := false;
    variable goto_L4341 : boolean := false;
    variable goto_L4338 : boolean := false;
    variable goto_L4382 : boolean := false;
    variable goto_L4393 : boolean := false;
    variable goto_L4404 : boolean := false;
    variable goto_L4396 : boolean := false;
    variable goto_L4385 : boolean := false;
    variable goto_L4374 : boolean := false;
    variable goto_L4371 : boolean := false;
    variable goto_L4138 : boolean := false;
    variable goto_L4051 : boolean := false;
    variable goto_L3990 : boolean := false;
    variable goto_L3895 : boolean := false;
    variable goto_L3908 : boolean := false;
    variable goto_L3915 : boolean := false;
    variable goto_L3922 : boolean := false;
    variable goto_L3918 : boolean := false;
    variable goto_L3911 : boolean := false;
    variable goto_L3904 : boolean := false;
    variable goto_L3901 : boolean := false;
    variable goto_L3784 : boolean := false;
    variable goto_L3836 : boolean := false;
    variable goto_L3795 : boolean := false;
    variable goto_L3808 : boolean := false;
    variable goto_L3815 : boolean := false;
    variable goto_L3822 : boolean := false;
    variable goto_L3818 : boolean := false;
    variable goto_L3811 : boolean := false;
    variable goto_L3804 : boolean := false;
    variable goto_L3801 : boolean := false;
    variable goto_L3791 : boolean := false;
    variable goto_L3675 : boolean := false;
    variable goto_L3725 : boolean := false;
    variable goto_L3684 : boolean := false;
    variable goto_L3697 : boolean := false;
    variable goto_L3704 : boolean := false;
    variable goto_L3711 : boolean := false;
    variable goto_L3707 : boolean := false;
    variable goto_L3700 : boolean := false;
    variable goto_L3693 : boolean := false;
    variable goto_L3690 : boolean := false;
    variable goto_L3680 : boolean := false;
    variable goto_L3564 : boolean := false;
    variable goto_L3616 : boolean := false;
    variable goto_L3575 : boolean := false;
    variable goto_L3588 : boolean := false;
    variable goto_L3595 : boolean := false;
    variable goto_L3602 : boolean := false;
    variable goto_L3598 : boolean := false;
    variable goto_L3591 : boolean := false;
    variable goto_L3584 : boolean := false;
    variable goto_L3581 : boolean := false;
    variable goto_L3571 : boolean := false;
    variable goto_L3455 : boolean := false;
    variable goto_L3505 : boolean := false;
    variable goto_L3464 : boolean := false;
    variable goto_L3477 : boolean := false;
    variable goto_L3484 : boolean := false;
    variable goto_L3491 : boolean := false;
    variable goto_L3487 : boolean := false;
    variable goto_L3480 : boolean := false;
    variable goto_L3473 : boolean := false;
    variable goto_L3470 : boolean := false;
    variable goto_L3460 : boolean := false;
    variable goto_L3281 : boolean := false;
    variable goto_L3294 : boolean := false;
    variable goto_L3301 : boolean := false;
    variable goto_L3308 : boolean := false;
    variable goto_L3304 : boolean := false;
    variable goto_L3297 : boolean := false;
    variable goto_L3290 : boolean := false;
    variable goto_L3287 : boolean := false;
    variable goto_L3328 : boolean := false;
    variable goto_L3335 : boolean := false;
    variable goto_L3342 : boolean := false;
    variable goto_L3338 : boolean := false;
    variable goto_L3331 : boolean := false;
    variable goto_L3324 : boolean := false;
    variable goto_L3321 : boolean := false;
    variable goto_L3095 : boolean := false;
    variable goto_L3108 : boolean := false;
    variable goto_L3115 : boolean := false;
    variable goto_L3122 : boolean := false;
    variable goto_L3118 : boolean := false;
    variable goto_L3111 : boolean := false;
    variable goto_L3104 : boolean := false;
    variable goto_L3101 : boolean := false;
    variable goto_L3142 : boolean := false;
    variable goto_L3149 : boolean := false;
    variable goto_L3156 : boolean := false;
    variable goto_L3152 : boolean := false;
    variable goto_L3145 : boolean := false;
    variable goto_L3138 : boolean := false;
    variable goto_L3135 : boolean := false;
    variable goto_L3181 : boolean := false;
    variable goto_L3190 : boolean := false;
    variable goto_L3199 : boolean := false;
    variable goto_L3193 : boolean := false;
    variable goto_L3184 : boolean := false;
    variable goto_L3175 : boolean := false;
    variable goto_L3172 : boolean := false;
    variable goto_L2909 : boolean := false;
    variable goto_L2922 : boolean := false;
    variable goto_L2929 : boolean := false;
    variable goto_L2936 : boolean := false;
    variable goto_L2932 : boolean := false;
    variable goto_L2925 : boolean := false;
    variable goto_L2918 : boolean := false;
    variable goto_L2915 : boolean := false;
    variable goto_L2956 : boolean := false;
    variable goto_L2963 : boolean := false;
    variable goto_L2970 : boolean := false;
    variable goto_L2966 : boolean := false;
    variable goto_L2959 : boolean := false;
    variable goto_L2952 : boolean := false;
    variable goto_L2949 : boolean := false;
    variable goto_L2995 : boolean := false;
    variable goto_L3004 : boolean := false;
    variable goto_L3013 : boolean := false;
    variable goto_L3007 : boolean := false;
    variable goto_L2998 : boolean := false;
    variable goto_L2989 : boolean := false;
    variable goto_L2986 : boolean := false;
    variable goto_L2723 : boolean := false;
    variable goto_L2736 : boolean := false;
    variable goto_L2743 : boolean := false;
    variable goto_L2750 : boolean := false;
    variable goto_L2746 : boolean := false;
    variable goto_L2739 : boolean := false;
    variable goto_L2732 : boolean := false;
    variable goto_L2729 : boolean := false;
    variable goto_L2770 : boolean := false;
    variable goto_L2777 : boolean := false;
    variable goto_L2784 : boolean := false;
    variable goto_L2780 : boolean := false;
    variable goto_L2773 : boolean := false;
    variable goto_L2766 : boolean := false;
    variable goto_L2763 : boolean := false;
    variable goto_L2809 : boolean := false;
    variable goto_L2818 : boolean := false;
    variable goto_L2827 : boolean := false;
    variable goto_L2821 : boolean := false;
    variable goto_L2812 : boolean := false;
    variable goto_L2803 : boolean := false;
    variable goto_L2800 : boolean := false;
    variable goto_L2594 : boolean := false;
    variable goto_L2607 : boolean := false;
    variable goto_L2614 : boolean := false;
    variable goto_L2621 : boolean := false;
    variable goto_L2617 : boolean := false;
    variable goto_L2610 : boolean := false;
    variable goto_L2603 : boolean := false;
    variable goto_L2600 : boolean := false;
    variable goto_L2642 : boolean := false;
    variable goto_L2651 : boolean := false;
    variable goto_L2660 : boolean := false;
    variable goto_L2654 : boolean := false;
    variable goto_L2645 : boolean := false;
    variable goto_L2636 : boolean := false;
    variable goto_L2633 : boolean := false;
    variable goto_L2386 : boolean := false;
    variable goto_L2399 : boolean := false;
    variable goto_L2406 : boolean := false;
    variable goto_L2413 : boolean := false;
    variable goto_L2409 : boolean := false;
    variable goto_L2402 : boolean := false;
    variable goto_L2395 : boolean := false;
    variable goto_L2392 : boolean := false;
    variable goto_L2433 : boolean := false;
    variable goto_L2440 : boolean := false;
    variable goto_L2447 : boolean := false;
    variable goto_L2443 : boolean := false;
    variable goto_L2436 : boolean := false;
    variable goto_L2429 : boolean := false;
    variable goto_L2426 : boolean := false;
    variable goto_L2513 : boolean := false;
    variable goto_L2522 : boolean := false;
    variable goto_L2531 : boolean := false;
    variable goto_L2525 : boolean := false;
    variable goto_L2516 : boolean := false;
    variable goto_L2507 : boolean := false;
    variable goto_L2504 : boolean := false;
    variable goto_L2182 : boolean := false;
    variable goto_L2195 : boolean := false;
    variable goto_L2202 : boolean := false;
    variable goto_L2209 : boolean := false;
    variable goto_L2205 : boolean := false;
    variable goto_L2198 : boolean := false;
    variable goto_L2191 : boolean := false;
    variable goto_L2188 : boolean := false;
    variable goto_L2229 : boolean := false;
    variable goto_L2236 : boolean := false;
    variable goto_L2243 : boolean := false;
    variable goto_L2239 : boolean := false;
    variable goto_L2232 : boolean := false;
    variable goto_L2225 : boolean := false;
    variable goto_L2222 : boolean := false;
    variable goto_L2305 : boolean := false;
    variable goto_L2314 : boolean := false;
    variable goto_L2323 : boolean := false;
    variable goto_L2317 : boolean := false;
    variable goto_L2308 : boolean := false;
    variable goto_L2299 : boolean := false;
    variable goto_L2296 : boolean := false;
    variable goto_L1974 : boolean := false;
    variable goto_L1987 : boolean := false;
    variable goto_L1994 : boolean := false;
    variable goto_L2001 : boolean := false;
    variable goto_L1997 : boolean := false;
    variable goto_L1990 : boolean := false;
    variable goto_L1983 : boolean := false;
    variable goto_L1980 : boolean := false;
    variable goto_L2021 : boolean := false;
    variable goto_L2028 : boolean := false;
    variable goto_L2035 : boolean := false;
    variable goto_L2031 : boolean := false;
    variable goto_L2024 : boolean := false;
    variable goto_L2017 : boolean := false;
    variable goto_L2014 : boolean := false;
    variable goto_L2101 : boolean := false;
    variable goto_L2110 : boolean := false;
    variable goto_L2119 : boolean := false;
    variable goto_L2113 : boolean := false;
    variable goto_L2104 : boolean := false;
    variable goto_L2095 : boolean := false;
    variable goto_L2092 : boolean := false;
    variable goto_L1770 : boolean := false;
    variable goto_L1783 : boolean := false;
    variable goto_L1790 : boolean := false;
    variable goto_L1797 : boolean := false;
    variable goto_L1793 : boolean := false;
    variable goto_L1786 : boolean := false;
    variable goto_L1779 : boolean := false;
    variable goto_L1776 : boolean := false;
    variable goto_L1817 : boolean := false;
    variable goto_L1824 : boolean := false;
    variable goto_L1831 : boolean := false;
    variable goto_L1827 : boolean := false;
    variable goto_L1820 : boolean := false;
    variable goto_L1813 : boolean := false;
    variable goto_L1810 : boolean := false;
    variable goto_L1893 : boolean := false;
    variable goto_L1902 : boolean := false;
    variable goto_L1911 : boolean := false;
    variable goto_L1905 : boolean := false;
    variable goto_L1896 : boolean := false;
    variable goto_L1887 : boolean := false;
    variable goto_L1884 : boolean := false;
    variable goto_L1602 : boolean := false;
    variable goto_L1615 : boolean := false;
    variable goto_L1622 : boolean := false;
    variable goto_L1629 : boolean := false;
    variable goto_L1625 : boolean := false;
    variable goto_L1618 : boolean := false;
    variable goto_L1611 : boolean := false;
    variable goto_L1608 : boolean := false;
    variable goto_L1649 : boolean := false;
    variable goto_L1656 : boolean := false;
    variable goto_L1663 : boolean := false;
    variable goto_L1659 : boolean := false;
    variable goto_L1652 : boolean := false;
    variable goto_L1645 : boolean := false;
    variable goto_L1642 : boolean := false;
    variable goto_L1434 : boolean := false;
    variable goto_L1447 : boolean := false;
    variable goto_L1454 : boolean := false;
    variable goto_L1461 : boolean := false;
    variable goto_L1457 : boolean := false;
    variable goto_L1450 : boolean := false;
    variable goto_L1443 : boolean := false;
    variable goto_L1440 : boolean := false;
    variable goto_L770 : boolean := false;
    variable goto_L418 : boolean := false;
    variable goto_L283 : boolean := false;
    variable goto_L0 : boolean := false;
    variable goto_L5439 : boolean := false;
    variable r5432 : std_logic_vector(0 to 80) := (others => '0');
    variable r5428 : std_logic_vector(0 to 80) := (others => '0');
    variable r5426 : std_logic_vector(0 to 9) := (others => '0');
    variable r5422 : std_logic_vector(0 to 17) := (others => '0');
    variable r5419 : std_logic_vector(0 to 80) := (others => '0');
    variable r5416 : std_logic_vector(0 to 80) := (others => '0');
    variable r5414 : std_logic_vector(0 to 17) := (others => '0');
    variable r5411 : std_logic_vector(0 to 80) := (others => '0');
    variable r5408 : std_logic_vector(0 to 80) := (others => '0');
    variable r5406 : std_logic_vector(0 to 0) := (others => '0');
    variable r5403 : std_logic_vector(0 to 80) := (others => '0');
    variable r5400 : std_logic_vector(0 to 80) := (others => '0');
    variable r5398 : std_logic_vector(0 to 0) := (others => '0');
    variable r5395 : std_logic_vector(0 to 80) := (others => '0');
    variable b5393 : boolean := false;
    variable r5388 : std_logic_vector(0 to 80) := (others => '0');
    variable r5384 : std_logic_vector(0 to 80) := (others => '0');
    variable r5382 : std_logic_vector(0 to 9) := (others => '0');
    variable r5378 : std_logic_vector(0 to 17) := (others => '0');
    variable r5375 : std_logic_vector(0 to 80) := (others => '0');
    variable r5372 : std_logic_vector(0 to 80) := (others => '0');
    variable r5370 : std_logic_vector(0 to 0) := (others => '0');
    variable r5368 : std_logic_vector(0 to 7) := (others => '0');
    variable r5364 : std_logic_vector(0 to 80) := (others => '0');
    variable r5361 : std_logic_vector(0 to 80) := (others => '0');
    variable r5357 : std_logic_vector(0 to 80) := (others => '0');
    variable r5353 : std_logic_vector(0 to 80) := (others => '0');
    variable r5345 : std_logic_vector(0 to 80) := (others => '0');
    variable b5341 : boolean := false;
    variable r5336 : std_logic_vector(0 to 80) := (others => '0');
    variable b5332 : boolean := false;
    variable r5327 : std_logic_vector(0 to 80) := (others => '0');
    variable b5323 : boolean := false;
    variable r5320 : std_logic_vector(0 to 1) := (others => '0');
    variable r5316 : std_logic_vector(0 to 80) := (others => '0');
    variable b5311 : boolean := false;
    variable b5309 : boolean := false;
    variable r5307 : std_logic_vector(0 to 7) := (others => '0');
    variable r5305 : std_logic_vector(0 to 0) := (others => '0');
    variable r5303 : std_logic_vector(0 to 7) := (others => '0');
    variable b5297 : boolean := false;
    variable b5295 : boolean := false;
    variable r5293 : std_logic_vector(0 to 7) := (others => '0');
    variable r5291 : std_logic_vector(0 to 0) := (others => '0');
    variable r5289 : std_logic_vector(0 to 0) := (others => '0');
    variable r5284 : std_logic_vector(0 to 8) := (others => '0');
    variable r5282 : std_logic_vector(0 to 0) := (others => '0');
    variable r5277 : std_logic_vector(0 to 0) := (others => '0');
    variable r5275 : std_logic_vector(0 to 0) := (others => '0');
    variable r5270 : std_logic_vector(0 to 8) := (others => '0');
    variable r5268 : std_logic_vector(0 to 0) := (others => '0');
    variable b5264 : boolean := false;
    variable b5262 : boolean := false;
    variable b5260 : boolean := false;
    variable r5258 : std_logic_vector(0 to 0) := (others => '0');
    variable r5256 : std_logic_vector(0 to 0) := (others => '0');
    variable b5254 : boolean := false;
    variable r5250 : std_logic_vector(0 to 8) := (others => '0');
    variable r5248 : std_logic_vector(0 to 0) := (others => '0');
    variable b5245 : boolean := false;
    variable b5243 : boolean := false;
    variable b5241 : boolean := false;
    variable r5239 : std_logic_vector(0 to 0) := (others => '0');
    variable r5237 : std_logic_vector(0 to 0) := (others => '0');
    variable b5235 : boolean := false;
    variable r5231 : std_logic_vector(0 to 8) := (others => '0');
    variable r5229 : std_logic_vector(0 to 0) := (others => '0');
    variable b5225 : boolean := false;
    variable b5223 : boolean := false;
    variable b5221 : boolean := false;
    variable r5219 : std_logic_vector(0 to 0) := (others => '0');
    variable r5217 : std_logic_vector(0 to 0) := (others => '0');
    variable b5215 : boolean := false;
    variable r5214 : std_logic_vector(0 to 8) := (others => '0');
    variable r5212 : std_logic_vector(0 to 1) := (others => '0');
    variable r5206 : std_logic_vector(0 to 7) := (others => '0');
    variable r5200 : std_logic_vector(0 to 7) := (others => '0');
    variable b5197 : boolean := false;
    variable r5193 : std_logic_vector(0 to 7) := (others => '0');
    variable b5190 : boolean := false;
    variable r5186 : std_logic_vector(0 to 7) := (others => '0');
    variable b5183 : boolean := false;
    variable r5181 : std_logic_vector(0 to 7) := (others => '0');
    variable r5179 : std_logic_vector(0 to 1) := (others => '0');
    variable r5175 : std_logic_vector(0 to 80) := (others => '0');
    variable b5173 : boolean := false;
    variable b5171 : boolean := false;
    variable b5169 : boolean := false;
    variable b5167 : boolean := false;
    variable b5165 : boolean := false;
    variable b5163 : boolean := false;
    variable b5161 : boolean := false;
    variable b5159 : boolean := false;
    variable b5157 : boolean := false;
    variable r5155 : std_logic_vector(0 to 0) := (others => '0');
    variable r5153 : std_logic_vector(0 to 0) := (others => '0');
    variable r5151 : std_logic_vector(0 to 0) := (others => '0');
    variable r5149 : std_logic_vector(0 to 0) := (others => '0');
    variable r5147 : std_logic_vector(0 to 0) := (others => '0');
    variable r5145 : std_logic_vector(0 to 0) := (others => '0');
    variable r5143 : std_logic_vector(0 to 0) := (others => '0');
    variable r5141 : std_logic_vector(0 to 0) := (others => '0');
    variable b5139 : boolean := false;
    variable r5133 : std_logic_vector(0 to 80) := (others => '0');
    variable r5129 : std_logic_vector(0 to 80) := (others => '0');
    variable r5127 : std_logic_vector(0 to 9) := (others => '0');
    variable r5123 : std_logic_vector(0 to 17) := (others => '0');
    variable r5120 : std_logic_vector(0 to 80) := (others => '0');
    variable r5116 : std_logic_vector(0 to 80) := (others => '0');
    variable r5114 : std_logic_vector(0 to 7) := (others => '0');
    variable r5106 : std_logic_vector(0 to 80) := (others => '0');
    variable r5104 : std_logic_vector(0 to 7) := (others => '0');
    variable b5100 : boolean := false;
    variable r5095 : std_logic_vector(0 to 80) := (others => '0');
    variable r5093 : std_logic_vector(0 to 7) := (others => '0');
    variable b5089 : boolean := false;
    variable r5084 : std_logic_vector(0 to 80) := (others => '0');
    variable r5082 : std_logic_vector(0 to 7) := (others => '0');
    variable b5078 : boolean := false;
    variable r5075 : std_logic_vector(0 to 1) := (others => '0');
    variable r5071 : std_logic_vector(0 to 80) := (others => '0');
    variable r5068 : std_logic_vector(0 to 7) := (others => '0');
    variable r5062 : std_logic_vector(0 to 7) := (others => '0');
    variable b5059 : boolean := false;
    variable r5055 : std_logic_vector(0 to 7) := (others => '0');
    variable b5052 : boolean := false;
    variable r5048 : std_logic_vector(0 to 7) := (others => '0');
    variable b5045 : boolean := false;
    variable r5043 : std_logic_vector(0 to 7) := (others => '0');
    variable r5041 : std_logic_vector(0 to 1) := (others => '0');
    variable r5037 : std_logic_vector(0 to 80) := (others => '0');
    variable r5031 : std_logic_vector(0 to 80) := (others => '0');
    variable r5027 : std_logic_vector(0 to 80) := (others => '0');
    variable r5025 : std_logic_vector(0 to 9) := (others => '0');
    variable r5021 : std_logic_vector(0 to 17) := (others => '0');
    variable r5018 : std_logic_vector(0 to 80) := (others => '0');
    variable r5014 : std_logic_vector(0 to 80) := (others => '0');
    variable r5012 : std_logic_vector(0 to 7) := (others => '0');
    variable r5004 : std_logic_vector(0 to 80) := (others => '0');
    variable r5002 : std_logic_vector(0 to 7) := (others => '0');
    variable b4998 : boolean := false;
    variable r4993 : std_logic_vector(0 to 80) := (others => '0');
    variable r4991 : std_logic_vector(0 to 7) := (others => '0');
    variable b4987 : boolean := false;
    variable r4982 : std_logic_vector(0 to 80) := (others => '0');
    variable r4980 : std_logic_vector(0 to 7) := (others => '0');
    variable b4976 : boolean := false;
    variable r4973 : std_logic_vector(0 to 1) := (others => '0');
    variable r4969 : std_logic_vector(0 to 80) := (others => '0');
    variable r4966 : std_logic_vector(0 to 7) := (others => '0');
    variable r4960 : std_logic_vector(0 to 7) := (others => '0');
    variable b4957 : boolean := false;
    variable r4953 : std_logic_vector(0 to 7) := (others => '0');
    variable b4950 : boolean := false;
    variable r4946 : std_logic_vector(0 to 7) := (others => '0');
    variable b4943 : boolean := false;
    variable r4941 : std_logic_vector(0 to 7) := (others => '0');
    variable r4939 : std_logic_vector(0 to 1) := (others => '0');
    variable r4935 : std_logic_vector(0 to 80) := (others => '0');
    variable b4933 : boolean := false;
    variable b4929 : boolean := false;
    variable b4927 : boolean := false;
    variable b4925 : boolean := false;
    variable b4923 : boolean := false;
    variable b4921 : boolean := false;
    variable b4919 : boolean := false;
    variable b4917 : boolean := false;
    variable b4915 : boolean := false;
    variable b4913 : boolean := false;
    variable r4911 : std_logic_vector(0 to 0) := (others => '0');
    variable r4909 : std_logic_vector(0 to 0) := (others => '0');
    variable r4907 : std_logic_vector(0 to 0) := (others => '0');
    variable r4905 : std_logic_vector(0 to 0) := (others => '0');
    variable r4903 : std_logic_vector(0 to 0) := (others => '0');
    variable r4901 : std_logic_vector(0 to 0) := (others => '0');
    variable r4899 : std_logic_vector(0 to 0) := (others => '0');
    variable r4897 : std_logic_vector(0 to 0) := (others => '0');
    variable b4895 : boolean := false;
    variable r4890 : std_logic_vector(0 to 80) := (others => '0');
    variable r4886 : std_logic_vector(0 to 80) := (others => '0');
    variable r4884 : std_logic_vector(0 to 9) := (others => '0');
    variable r4880 : std_logic_vector(0 to 17) := (others => '0');
    variable r4877 : std_logic_vector(0 to 80) := (others => '0');
    variable r4874 : std_logic_vector(0 to 80) := (others => '0');
    variable r4872 : std_logic_vector(0 to 0) := (others => '0');
    variable r4870 : std_logic_vector(0 to 7) := (others => '0');
    variable r4866 : std_logic_vector(0 to 80) := (others => '0');
    variable r4863 : std_logic_vector(0 to 80) := (others => '0');
    variable r4859 : std_logic_vector(0 to 80) := (others => '0');
    variable r4855 : std_logic_vector(0 to 80) := (others => '0');
    variable r4847 : std_logic_vector(0 to 80) := (others => '0');
    variable b4843 : boolean := false;
    variable r4838 : std_logic_vector(0 to 80) := (others => '0');
    variable b4834 : boolean := false;
    variable r4829 : std_logic_vector(0 to 80) := (others => '0');
    variable b4825 : boolean := false;
    variable r4822 : std_logic_vector(0 to 1) := (others => '0');
    variable r4818 : std_logic_vector(0 to 80) := (others => '0');
    variable b4813 : boolean := false;
    variable b4811 : boolean := false;
    variable r4809 : std_logic_vector(0 to 7) := (others => '0');
    variable r4807 : std_logic_vector(0 to 0) := (others => '0');
    variable r4805 : std_logic_vector(0 to 7) := (others => '0');
    variable b4799 : boolean := false;
    variable b4797 : boolean := false;
    variable r4795 : std_logic_vector(0 to 7) := (others => '0');
    variable r4793 : std_logic_vector(0 to 0) := (others => '0');
    variable r4791 : std_logic_vector(0 to 0) := (others => '0');
    variable r4788 : std_logic_vector(0 to 8) := (others => '0');
    variable r4786 : std_logic_vector(0 to 0) := (others => '0');
    variable r4784 : std_logic_vector(0 to 7) := (others => '0');
    variable r4780 : std_logic_vector(0 to 7) := (others => '0');
    variable r4774 : std_logic_vector(0 to 7) := (others => '0');
    variable b4771 : boolean := false;
    variable r4767 : std_logic_vector(0 to 7) := (others => '0');
    variable b4764 : boolean := false;
    variable r4760 : std_logic_vector(0 to 7) := (others => '0');
    variable b4757 : boolean := false;
    variable r4755 : std_logic_vector(0 to 7) := (others => '0');
    variable r4753 : std_logic_vector(0 to 1) := (others => '0');
    variable r4749 : std_logic_vector(0 to 80) := (others => '0');
    variable b4747 : boolean := false;
    variable b4745 : boolean := false;
    variable b4743 : boolean := false;
    variable b4741 : boolean := false;
    variable b4739 : boolean := false;
    variable b4737 : boolean := false;
    variable b4735 : boolean := false;
    variable b4733 : boolean := false;
    variable b4731 : boolean := false;
    variable r4729 : std_logic_vector(0 to 0) := (others => '0');
    variable r4727 : std_logic_vector(0 to 0) := (others => '0');
    variable r4725 : std_logic_vector(0 to 0) := (others => '0');
    variable r4723 : std_logic_vector(0 to 0) := (others => '0');
    variable r4721 : std_logic_vector(0 to 0) := (others => '0');
    variable r4719 : std_logic_vector(0 to 0) := (others => '0');
    variable r4717 : std_logic_vector(0 to 0) := (others => '0');
    variable r4715 : std_logic_vector(0 to 0) := (others => '0');
    variable b4713 : boolean := false;
    variable r4708 : std_logic_vector(0 to 80) := (others => '0');
    variable r4704 : std_logic_vector(0 to 80) := (others => '0');
    variable r4702 : std_logic_vector(0 to 9) := (others => '0');
    variable r4698 : std_logic_vector(0 to 17) := (others => '0');
    variable r4695 : std_logic_vector(0 to 80) := (others => '0');
    variable r4692 : std_logic_vector(0 to 80) := (others => '0');
    variable r4690 : std_logic_vector(0 to 0) := (others => '0');
    variable r4688 : std_logic_vector(0 to 7) := (others => '0');
    variable r4684 : std_logic_vector(0 to 80) := (others => '0');
    variable r4681 : std_logic_vector(0 to 80) := (others => '0');
    variable r4677 : std_logic_vector(0 to 80) := (others => '0');
    variable r4673 : std_logic_vector(0 to 80) := (others => '0');
    variable r4665 : std_logic_vector(0 to 80) := (others => '0');
    variable b4661 : boolean := false;
    variable r4656 : std_logic_vector(0 to 80) := (others => '0');
    variable b4652 : boolean := false;
    variable r4647 : std_logic_vector(0 to 80) := (others => '0');
    variable b4643 : boolean := false;
    variable r4640 : std_logic_vector(0 to 1) := (others => '0');
    variable r4636 : std_logic_vector(0 to 80) := (others => '0');
    variable b4631 : boolean := false;
    variable b4629 : boolean := false;
    variable r4627 : std_logic_vector(0 to 7) := (others => '0');
    variable r4625 : std_logic_vector(0 to 0) := (others => '0');
    variable r4623 : std_logic_vector(0 to 7) := (others => '0');
    variable b4617 : boolean := false;
    variable b4615 : boolean := false;
    variable r4613 : std_logic_vector(0 to 7) := (others => '0');
    variable r4611 : std_logic_vector(0 to 0) := (others => '0');
    variable r4609 : std_logic_vector(0 to 0) := (others => '0');
    variable r4606 : std_logic_vector(0 to 8) := (others => '0');
    variable r4604 : std_logic_vector(0 to 0) := (others => '0');
    variable r4602 : std_logic_vector(0 to 7) := (others => '0');
    variable r4598 : std_logic_vector(0 to 7) := (others => '0');
    variable r4592 : std_logic_vector(0 to 7) := (others => '0');
    variable b4589 : boolean := false;
    variable r4585 : std_logic_vector(0 to 7) := (others => '0');
    variable b4582 : boolean := false;
    variable r4578 : std_logic_vector(0 to 7) := (others => '0');
    variable b4575 : boolean := false;
    variable r4573 : std_logic_vector(0 to 7) := (others => '0');
    variable r4571 : std_logic_vector(0 to 1) := (others => '0');
    variable r4567 : std_logic_vector(0 to 80) := (others => '0');
    variable b4565 : boolean := false;
    variable b4563 : boolean := false;
    variable b4561 : boolean := false;
    variable b4559 : boolean := false;
    variable b4557 : boolean := false;
    variable b4555 : boolean := false;
    variable b4553 : boolean := false;
    variable b4551 : boolean := false;
    variable b4549 : boolean := false;
    variable r4547 : std_logic_vector(0 to 0) := (others => '0');
    variable r4545 : std_logic_vector(0 to 0) := (others => '0');
    variable r4543 : std_logic_vector(0 to 0) := (others => '0');
    variable r4541 : std_logic_vector(0 to 0) := (others => '0');
    variable r4539 : std_logic_vector(0 to 0) := (others => '0');
    variable r4537 : std_logic_vector(0 to 0) := (others => '0');
    variable r4535 : std_logic_vector(0 to 0) := (others => '0');
    variable r4533 : std_logic_vector(0 to 0) := (others => '0');
    variable b4531 : boolean := false;
    variable r4526 : std_logic_vector(0 to 80) := (others => '0');
    variable r4522 : std_logic_vector(0 to 80) := (others => '0');
    variable r4520 : std_logic_vector(0 to 9) := (others => '0');
    variable r4516 : std_logic_vector(0 to 17) := (others => '0');
    variable r4513 : std_logic_vector(0 to 80) := (others => '0');
    variable r4509 : std_logic_vector(0 to 80) := (others => '0');
    variable r4507 : std_logic_vector(0 to 7) := (others => '0');
    variable r4500 : std_logic_vector(0 to 80) := (others => '0');
    variable r4498 : std_logic_vector(0 to 7) := (others => '0');
    variable b4495 : boolean := false;
    variable r4490 : std_logic_vector(0 to 80) := (others => '0');
    variable r4488 : std_logic_vector(0 to 7) := (others => '0');
    variable b4485 : boolean := false;
    variable r4480 : std_logic_vector(0 to 80) := (others => '0');
    variable r4478 : std_logic_vector(0 to 7) := (others => '0');
    variable b4475 : boolean := false;
    variable r4472 : std_logic_vector(0 to 1) := (others => '0');
    variable r4468 : std_logic_vector(0 to 80) := (others => '0');
    variable b4466 : boolean := false;
    variable b4464 : boolean := false;
    variable b4462 : boolean := false;
    variable b4460 : boolean := false;
    variable b4458 : boolean := false;
    variable b4456 : boolean := false;
    variable b4454 : boolean := false;
    variable b4452 : boolean := false;
    variable b4450 : boolean := false;
    variable r4448 : std_logic_vector(0 to 0) := (others => '0');
    variable r4446 : std_logic_vector(0 to 0) := (others => '0');
    variable r4444 : std_logic_vector(0 to 0) := (others => '0');
    variable r4442 : std_logic_vector(0 to 0) := (others => '0');
    variable r4440 : std_logic_vector(0 to 0) := (others => '0');
    variable r4438 : std_logic_vector(0 to 0) := (others => '0');
    variable r4436 : std_logic_vector(0 to 0) := (others => '0');
    variable r4434 : std_logic_vector(0 to 0) := (others => '0');
    variable b4432 : boolean := false;
    variable r4427 : std_logic_vector(0 to 80) := (others => '0');
    variable r4423 : std_logic_vector(0 to 80) := (others => '0');
    variable r4421 : std_logic_vector(0 to 9) := (others => '0');
    variable r4417 : std_logic_vector(0 to 17) := (others => '0');
    variable r4414 : std_logic_vector(0 to 80) := (others => '0');
    variable r4410 : std_logic_vector(0 to 80) := (others => '0');
    variable r4408 : std_logic_vector(0 to 7) := (others => '0');
    variable r4400 : std_logic_vector(0 to 80) := (others => '0');
    variable r4398 : std_logic_vector(0 to 7) := (others => '0');
    variable b4394 : boolean := false;
    variable r4389 : std_logic_vector(0 to 80) := (others => '0');
    variable r4387 : std_logic_vector(0 to 7) := (others => '0');
    variable b4383 : boolean := false;
    variable r4378 : std_logic_vector(0 to 80) := (others => '0');
    variable r4376 : std_logic_vector(0 to 7) := (others => '0');
    variable b4372 : boolean := false;
    variable r4369 : std_logic_vector(0 to 1) := (others => '0');
    variable r4365 : std_logic_vector(0 to 80) := (others => '0');
    variable r4362 : std_logic_vector(0 to 7) := (others => '0');
    variable r4356 : std_logic_vector(0 to 7) := (others => '0');
    variable b4353 : boolean := false;
    variable r4349 : std_logic_vector(0 to 7) := (others => '0');
    variable b4346 : boolean := false;
    variable r4342 : std_logic_vector(0 to 7) := (others => '0');
    variable b4339 : boolean := false;
    variable r4337 : std_logic_vector(0 to 7) := (others => '0');
    variable r4335 : std_logic_vector(0 to 1) := (others => '0');
    variable r4331 : std_logic_vector(0 to 80) := (others => '0');
    variable b4329 : boolean := false;
    variable b4327 : boolean := false;
    variable b4325 : boolean := false;
    variable b4323 : boolean := false;
    variable b4321 : boolean := false;
    variable b4319 : boolean := false;
    variable b4317 : boolean := false;
    variable b4315 : boolean := false;
    variable b4313 : boolean := false;
    variable r4311 : std_logic_vector(0 to 0) := (others => '0');
    variable r4309 : std_logic_vector(0 to 0) := (others => '0');
    variable r4307 : std_logic_vector(0 to 0) := (others => '0');
    variable r4305 : std_logic_vector(0 to 0) := (others => '0');
    variable r4303 : std_logic_vector(0 to 0) := (others => '0');
    variable r4301 : std_logic_vector(0 to 0) := (others => '0');
    variable r4299 : std_logic_vector(0 to 0) := (others => '0');
    variable r4297 : std_logic_vector(0 to 0) := (others => '0');
    variable b4295 : boolean := false;
    variable r4290 : std_logic_vector(0 to 80) := (others => '0');
    variable r4286 : std_logic_vector(0 to 80) := (others => '0');
    variable r4284 : std_logic_vector(0 to 9) := (others => '0');
    variable r4280 : std_logic_vector(0 to 17) := (others => '0');
    variable r4277 : std_logic_vector(0 to 80) := (others => '0');
    variable r4274 : std_logic_vector(0 to 80) := (others => '0');
    variable r4270 : std_logic_vector(0 to 80) := (others => '0');
    variable r4268 : std_logic_vector(0 to 0) := (others => '0');
    variable r4237 : std_logic_vector(0 to 0) := (others => '0');
    variable r4236 : std_logic_vector(0 to 80) := (others => '0');
    variable r4233 : std_logic_vector(0 to 80) := (others => '0');
    variable r4230 : std_logic_vector(0 to 80) := (others => '0');
    variable r4226 : std_logic_vector(0 to 80) := (others => '0');
    variable r4224 : std_logic_vector(0 to 0) := (others => '0');
    variable r4193 : std_logic_vector(0 to 0) := (others => '0');
    variable r4192 : std_logic_vector(0 to 80) := (others => '0');
    variable r4189 : std_logic_vector(0 to 80) := (others => '0');
    variable r4186 : std_logic_vector(0 to 80) := (others => '0');
    variable r4182 : std_logic_vector(0 to 80) := (others => '0');
    variable r4180 : std_logic_vector(0 to 7) := (others => '0');
    variable r4149 : std_logic_vector(0 to 7) := (others => '0');
    variable r4148 : std_logic_vector(0 to 80) := (others => '0');
    variable r4145 : std_logic_vector(0 to 80) := (others => '0');
    variable r4142 : std_logic_vector(0 to 80) := (others => '0');
    variable r4140 : std_logic_vector(0 to 0) := (others => '0');
    variable r4137 : std_logic_vector(0 to 80) := (others => '0');
    variable b4135 : boolean := false;
    variable b4133 : boolean := false;
    variable b4131 : boolean := false;
    variable b4129 : boolean := false;
    variable b4127 : boolean := false;
    variable b4125 : boolean := false;
    variable b4123 : boolean := false;
    variable b4121 : boolean := false;
    variable b4119 : boolean := false;
    variable r4117 : std_logic_vector(0 to 0) := (others => '0');
    variable r4115 : std_logic_vector(0 to 0) := (others => '0');
    variable r4113 : std_logic_vector(0 to 0) := (others => '0');
    variable r4111 : std_logic_vector(0 to 0) := (others => '0');
    variable r4109 : std_logic_vector(0 to 0) := (others => '0');
    variable r4107 : std_logic_vector(0 to 0) := (others => '0');
    variable r4105 : std_logic_vector(0 to 0) := (others => '0');
    variable r4103 : std_logic_vector(0 to 0) := (others => '0');
    variable b4101 : boolean := false;
    variable r4096 : std_logic_vector(0 to 80) := (others => '0');
    variable r4092 : std_logic_vector(0 to 80) := (others => '0');
    variable r4090 : std_logic_vector(0 to 9) := (others => '0');
    variable r4086 : std_logic_vector(0 to 17) := (others => '0');
    variable r4083 : std_logic_vector(0 to 80) := (others => '0');
    variable r4080 : std_logic_vector(0 to 80) := (others => '0');
    variable r4078 : std_logic_vector(0 to 17) := (others => '0');
    variable r4076 : std_logic_vector(0 to 0) := (others => '0');
    variable r4061 : std_logic_vector(0 to 17) := (others => '0');
    variable r4060 : std_logic_vector(0 to 0) := (others => '0');
    variable r4059 : std_logic_vector(0 to 17) := (others => '0');
    variable r4055 : std_logic_vector(0 to 80) := (others => '0');
    variable r4053 : std_logic_vector(0 to 17) := (others => '0');
    variable r4050 : std_logic_vector(0 to 80) := (others => '0');
    variable b4048 : boolean := false;
    variable b4046 : boolean := false;
    variable b4044 : boolean := false;
    variable b4042 : boolean := false;
    variable b4040 : boolean := false;
    variable b4038 : boolean := false;
    variable b4036 : boolean := false;
    variable b4034 : boolean := false;
    variable b4032 : boolean := false;
    variable r4030 : std_logic_vector(0 to 0) := (others => '0');
    variable r4028 : std_logic_vector(0 to 0) := (others => '0');
    variable r4026 : std_logic_vector(0 to 0) := (others => '0');
    variable r4024 : std_logic_vector(0 to 0) := (others => '0');
    variable r4022 : std_logic_vector(0 to 0) := (others => '0');
    variable r4020 : std_logic_vector(0 to 0) := (others => '0');
    variable r4018 : std_logic_vector(0 to 0) := (others => '0');
    variable r4016 : std_logic_vector(0 to 0) := (others => '0');
    variable b4014 : boolean := false;
    variable r4009 : std_logic_vector(0 to 80) := (others => '0');
    variable r4005 : std_logic_vector(0 to 80) := (others => '0');
    variable r4003 : std_logic_vector(0 to 9) := (others => '0');
    variable r3999 : std_logic_vector(0 to 17) := (others => '0');
    variable r3996 : std_logic_vector(0 to 80) := (others => '0');
    variable r3993 : std_logic_vector(0 to 80) := (others => '0');
    variable r3989 : std_logic_vector(0 to 80) := (others => '0');
    variable b3987 : boolean := false;
    variable b3985 : boolean := false;
    variable b3983 : boolean := false;
    variable b3981 : boolean := false;
    variable b3979 : boolean := false;
    variable b3977 : boolean := false;
    variable b3975 : boolean := false;
    variable b3973 : boolean := false;
    variable b3971 : boolean := false;
    variable r3969 : std_logic_vector(0 to 0) := (others => '0');
    variable r3967 : std_logic_vector(0 to 0) := (others => '0');
    variable r3965 : std_logic_vector(0 to 0) := (others => '0');
    variable r3963 : std_logic_vector(0 to 0) := (others => '0');
    variable r3961 : std_logic_vector(0 to 0) := (others => '0');
    variable r3959 : std_logic_vector(0 to 0) := (others => '0');
    variable r3957 : std_logic_vector(0 to 0) := (others => '0');
    variable r3955 : std_logic_vector(0 to 0) := (others => '0');
    variable b3953 : boolean := false;
    variable r3948 : std_logic_vector(0 to 80) := (others => '0');
    variable r3944 : std_logic_vector(0 to 80) := (others => '0');
    variable r3942 : std_logic_vector(0 to 9) := (others => '0');
    variable r3938 : std_logic_vector(0 to 17) := (others => '0');
    variable r3935 : std_logic_vector(0 to 80) := (others => '0');
    variable r3932 : std_logic_vector(0 to 80) := (others => '0');
    variable r3928 : std_logic_vector(0 to 80) := (others => '0');
    variable r3925 : std_logic_vector(0 to 7) := (others => '0');
    variable r3919 : std_logic_vector(0 to 7) := (others => '0');
    variable b3916 : boolean := false;
    variable r3912 : std_logic_vector(0 to 7) := (others => '0');
    variable b3909 : boolean := false;
    variable r3905 : std_logic_vector(0 to 7) := (others => '0');
    variable b3902 : boolean := false;
    variable r3900 : std_logic_vector(0 to 7) := (others => '0');
    variable r3898 : std_logic_vector(0 to 1) := (others => '0');
    variable r3894 : std_logic_vector(0 to 80) := (others => '0');
    variable b3892 : boolean := false;
    variable b3890 : boolean := false;
    variable b3888 : boolean := false;
    variable b3886 : boolean := false;
    variable b3884 : boolean := false;
    variable b3882 : boolean := false;
    variable b3880 : boolean := false;
    variable b3878 : boolean := false;
    variable b3876 : boolean := false;
    variable r3874 : std_logic_vector(0 to 0) := (others => '0');
    variable r3872 : std_logic_vector(0 to 0) := (others => '0');
    variable r3870 : std_logic_vector(0 to 0) := (others => '0');
    variable r3868 : std_logic_vector(0 to 0) := (others => '0');
    variable r3866 : std_logic_vector(0 to 0) := (others => '0');
    variable r3864 : std_logic_vector(0 to 0) := (others => '0');
    variable r3862 : std_logic_vector(0 to 0) := (others => '0');
    variable r3860 : std_logic_vector(0 to 0) := (others => '0');
    variable b3858 : boolean := false;
    variable r3853 : std_logic_vector(0 to 80) := (others => '0');
    variable r3849 : std_logic_vector(0 to 80) := (others => '0');
    variable r3847 : std_logic_vector(0 to 9) := (others => '0');
    variable r3843 : std_logic_vector(0 to 17) := (others => '0');
    variable r3840 : std_logic_vector(0 to 80) := (others => '0');
    variable r3832 : std_logic_vector(0 to 80) := (others => '0');
    variable r3828 : std_logic_vector(0 to 80) := (others => '0');
    variable r3825 : std_logic_vector(0 to 7) := (others => '0');
    variable r3819 : std_logic_vector(0 to 7) := (others => '0');
    variable b3816 : boolean := false;
    variable r3812 : std_logic_vector(0 to 7) := (others => '0');
    variable b3809 : boolean := false;
    variable r3805 : std_logic_vector(0 to 7) := (others => '0');
    variable b3802 : boolean := false;
    variable r3800 : std_logic_vector(0 to 7) := (others => '0');
    variable r3798 : std_logic_vector(0 to 1) := (others => '0');
    variable r3794 : std_logic_vector(0 to 80) := (others => '0');
    variable b3792 : boolean := false;
    variable r3789 : std_logic_vector(0 to 0) := (others => '0');
    variable r3786 : std_logic_vector(0 to 0) := (others => '0');
    variable r3783 : std_logic_vector(0 to 80) := (others => '0');
    variable b3781 : boolean := false;
    variable b3779 : boolean := false;
    variable b3777 : boolean := false;
    variable b3775 : boolean := false;
    variable b3773 : boolean := false;
    variable b3771 : boolean := false;
    variable b3769 : boolean := false;
    variable b3767 : boolean := false;
    variable b3765 : boolean := false;
    variable r3763 : std_logic_vector(0 to 0) := (others => '0');
    variable r3761 : std_logic_vector(0 to 0) := (others => '0');
    variable r3759 : std_logic_vector(0 to 0) := (others => '0');
    variable r3757 : std_logic_vector(0 to 0) := (others => '0');
    variable r3755 : std_logic_vector(0 to 0) := (others => '0');
    variable r3753 : std_logic_vector(0 to 0) := (others => '0');
    variable r3751 : std_logic_vector(0 to 0) := (others => '0');
    variable r3749 : std_logic_vector(0 to 0) := (others => '0');
    variable b3747 : boolean := false;
    variable r3742 : std_logic_vector(0 to 80) := (others => '0');
    variable r3738 : std_logic_vector(0 to 80) := (others => '0');
    variable r3736 : std_logic_vector(0 to 9) := (others => '0');
    variable r3732 : std_logic_vector(0 to 17) := (others => '0');
    variable r3729 : std_logic_vector(0 to 80) := (others => '0');
    variable r3721 : std_logic_vector(0 to 80) := (others => '0');
    variable r3717 : std_logic_vector(0 to 80) := (others => '0');
    variable r3714 : std_logic_vector(0 to 7) := (others => '0');
    variable r3708 : std_logic_vector(0 to 7) := (others => '0');
    variable b3705 : boolean := false;
    variable r3701 : std_logic_vector(0 to 7) := (others => '0');
    variable b3698 : boolean := false;
    variable r3694 : std_logic_vector(0 to 7) := (others => '0');
    variable b3691 : boolean := false;
    variable r3689 : std_logic_vector(0 to 7) := (others => '0');
    variable r3687 : std_logic_vector(0 to 1) := (others => '0');
    variable r3683 : std_logic_vector(0 to 80) := (others => '0');
    variable b3681 : boolean := false;
    variable r3677 : std_logic_vector(0 to 0) := (others => '0');
    variable r3674 : std_logic_vector(0 to 80) := (others => '0');
    variable b3672 : boolean := false;
    variable b3670 : boolean := false;
    variable b3668 : boolean := false;
    variable b3666 : boolean := false;
    variable b3664 : boolean := false;
    variable b3662 : boolean := false;
    variable b3660 : boolean := false;
    variable b3658 : boolean := false;
    variable b3656 : boolean := false;
    variable r3654 : std_logic_vector(0 to 0) := (others => '0');
    variable r3652 : std_logic_vector(0 to 0) := (others => '0');
    variable r3650 : std_logic_vector(0 to 0) := (others => '0');
    variable r3648 : std_logic_vector(0 to 0) := (others => '0');
    variable r3646 : std_logic_vector(0 to 0) := (others => '0');
    variable r3644 : std_logic_vector(0 to 0) := (others => '0');
    variable r3642 : std_logic_vector(0 to 0) := (others => '0');
    variable r3640 : std_logic_vector(0 to 0) := (others => '0');
    variable b3638 : boolean := false;
    variable r3633 : std_logic_vector(0 to 80) := (others => '0');
    variable r3629 : std_logic_vector(0 to 80) := (others => '0');
    variable r3627 : std_logic_vector(0 to 9) := (others => '0');
    variable r3623 : std_logic_vector(0 to 17) := (others => '0');
    variable r3620 : std_logic_vector(0 to 80) := (others => '0');
    variable r3612 : std_logic_vector(0 to 80) := (others => '0');
    variable r3608 : std_logic_vector(0 to 80) := (others => '0');
    variable r3605 : std_logic_vector(0 to 7) := (others => '0');
    variable r3599 : std_logic_vector(0 to 7) := (others => '0');
    variable b3596 : boolean := false;
    variable r3592 : std_logic_vector(0 to 7) := (others => '0');
    variable b3589 : boolean := false;
    variable r3585 : std_logic_vector(0 to 7) := (others => '0');
    variable b3582 : boolean := false;
    variable r3580 : std_logic_vector(0 to 7) := (others => '0');
    variable r3578 : std_logic_vector(0 to 1) := (others => '0');
    variable r3574 : std_logic_vector(0 to 80) := (others => '0');
    variable b3572 : boolean := false;
    variable r3569 : std_logic_vector(0 to 0) := (others => '0');
    variable r3566 : std_logic_vector(0 to 0) := (others => '0');
    variable r3563 : std_logic_vector(0 to 80) := (others => '0');
    variable b3561 : boolean := false;
    variable b3559 : boolean := false;
    variable b3557 : boolean := false;
    variable b3555 : boolean := false;
    variable b3553 : boolean := false;
    variable b3551 : boolean := false;
    variable b3549 : boolean := false;
    variable b3547 : boolean := false;
    variable b3545 : boolean := false;
    variable r3543 : std_logic_vector(0 to 0) := (others => '0');
    variable r3541 : std_logic_vector(0 to 0) := (others => '0');
    variable r3539 : std_logic_vector(0 to 0) := (others => '0');
    variable r3537 : std_logic_vector(0 to 0) := (others => '0');
    variable r3535 : std_logic_vector(0 to 0) := (others => '0');
    variable r3533 : std_logic_vector(0 to 0) := (others => '0');
    variable r3531 : std_logic_vector(0 to 0) := (others => '0');
    variable r3529 : std_logic_vector(0 to 0) := (others => '0');
    variable b3527 : boolean := false;
    variable r3522 : std_logic_vector(0 to 80) := (others => '0');
    variable r3518 : std_logic_vector(0 to 80) := (others => '0');
    variable r3516 : std_logic_vector(0 to 9) := (others => '0');
    variable r3512 : std_logic_vector(0 to 17) := (others => '0');
    variable r3509 : std_logic_vector(0 to 80) := (others => '0');
    variable r3501 : std_logic_vector(0 to 80) := (others => '0');
    variable r3497 : std_logic_vector(0 to 80) := (others => '0');
    variable r3494 : std_logic_vector(0 to 7) := (others => '0');
    variable r3488 : std_logic_vector(0 to 7) := (others => '0');
    variable b3485 : boolean := false;
    variable r3481 : std_logic_vector(0 to 7) := (others => '0');
    variable b3478 : boolean := false;
    variable r3474 : std_logic_vector(0 to 7) := (others => '0');
    variable b3471 : boolean := false;
    variable r3469 : std_logic_vector(0 to 7) := (others => '0');
    variable r3467 : std_logic_vector(0 to 1) := (others => '0');
    variable r3463 : std_logic_vector(0 to 80) := (others => '0');
    variable b3461 : boolean := false;
    variable r3457 : std_logic_vector(0 to 0) := (others => '0');
    variable r3454 : std_logic_vector(0 to 80) := (others => '0');
    variable b3452 : boolean := false;
    variable b3450 : boolean := false;
    variable b3448 : boolean := false;
    variable b3446 : boolean := false;
    variable b3444 : boolean := false;
    variable b3442 : boolean := false;
    variable b3440 : boolean := false;
    variable b3438 : boolean := false;
    variable b3436 : boolean := false;
    variable r3434 : std_logic_vector(0 to 0) := (others => '0');
    variable r3432 : std_logic_vector(0 to 0) := (others => '0');
    variable r3430 : std_logic_vector(0 to 0) := (others => '0');
    variable r3428 : std_logic_vector(0 to 0) := (others => '0');
    variable r3426 : std_logic_vector(0 to 0) := (others => '0');
    variable r3424 : std_logic_vector(0 to 0) := (others => '0');
    variable r3422 : std_logic_vector(0 to 0) := (others => '0');
    variable r3420 : std_logic_vector(0 to 0) := (others => '0');
    variable b3418 : boolean := false;
    variable r3413 : std_logic_vector(0 to 80) := (others => '0');
    variable r3409 : std_logic_vector(0 to 80) := (others => '0');
    variable r3407 : std_logic_vector(0 to 9) := (others => '0');
    variable r3403 : std_logic_vector(0 to 17) := (others => '0');
    variable r3400 : std_logic_vector(0 to 80) := (others => '0');
    variable r3397 : std_logic_vector(0 to 80) := (others => '0');
    variable r3395 : std_logic_vector(0 to 0) := (others => '0');
    variable r3393 : std_logic_vector(0 to 7) := (others => '0');
    variable r3389 : std_logic_vector(0 to 80) := (others => '0');
    variable r3386 : std_logic_vector(0 to 80) := (others => '0');
    variable r3382 : std_logic_vector(0 to 80) := (others => '0');
    variable b3377 : boolean := false;
    variable b3375 : boolean := false;
    variable r3373 : std_logic_vector(0 to 7) := (others => '0');
    variable r3371 : std_logic_vector(0 to 0) := (others => '0');
    variable r3369 : std_logic_vector(0 to 7) := (others => '0');
    variable b3363 : boolean := false;
    variable b3361 : boolean := false;
    variable r3359 : std_logic_vector(0 to 7) := (others => '0');
    variable r3357 : std_logic_vector(0 to 0) := (others => '0');
    variable r3355 : std_logic_vector(0 to 0) := (others => '0');
    variable r3352 : std_logic_vector(0 to 8) := (others => '0');
    variable r3350 : std_logic_vector(0 to 0) := (others => '0');
    variable r3345 : std_logic_vector(0 to 7) := (others => '0');
    variable r3339 : std_logic_vector(0 to 7) := (others => '0');
    variable b3336 : boolean := false;
    variable r3332 : std_logic_vector(0 to 7) := (others => '0');
    variable b3329 : boolean := false;
    variable r3325 : std_logic_vector(0 to 7) := (others => '0');
    variable b3322 : boolean := false;
    variable r3320 : std_logic_vector(0 to 7) := (others => '0');
    variable r3318 : std_logic_vector(0 to 1) := (others => '0');
    variable r3314 : std_logic_vector(0 to 80) := (others => '0');
    variable r3311 : std_logic_vector(0 to 7) := (others => '0');
    variable r3305 : std_logic_vector(0 to 7) := (others => '0');
    variable b3302 : boolean := false;
    variable r3298 : std_logic_vector(0 to 7) := (others => '0');
    variable b3295 : boolean := false;
    variable r3291 : std_logic_vector(0 to 7) := (others => '0');
    variable b3288 : boolean := false;
    variable r3286 : std_logic_vector(0 to 7) := (others => '0');
    variable r3284 : std_logic_vector(0 to 1) := (others => '0');
    variable r3280 : std_logic_vector(0 to 80) := (others => '0');
    variable b3278 : boolean := false;
    variable b3276 : boolean := false;
    variable b3274 : boolean := false;
    variable b3272 : boolean := false;
    variable b3270 : boolean := false;
    variable b3268 : boolean := false;
    variable b3266 : boolean := false;
    variable b3264 : boolean := false;
    variable b3262 : boolean := false;
    variable r3260 : std_logic_vector(0 to 0) := (others => '0');
    variable r3258 : std_logic_vector(0 to 0) := (others => '0');
    variable r3256 : std_logic_vector(0 to 0) := (others => '0');
    variable r3254 : std_logic_vector(0 to 0) := (others => '0');
    variable r3252 : std_logic_vector(0 to 0) := (others => '0');
    variable r3250 : std_logic_vector(0 to 0) := (others => '0');
    variable r3248 : std_logic_vector(0 to 0) := (others => '0');
    variable r3246 : std_logic_vector(0 to 0) := (others => '0');
    variable b3244 : boolean := false;
    variable r3239 : std_logic_vector(0 to 80) := (others => '0');
    variable r3235 : std_logic_vector(0 to 80) := (others => '0');
    variable r3233 : std_logic_vector(0 to 9) := (others => '0');
    variable r3229 : std_logic_vector(0 to 17) := (others => '0');
    variable r3226 : std_logic_vector(0 to 80) := (others => '0');
    variable r3223 : std_logic_vector(0 to 80) := (others => '0');
    variable r3221 : std_logic_vector(0 to 0) := (others => '0');
    variable r3219 : std_logic_vector(0 to 7) := (others => '0');
    variable r3215 : std_logic_vector(0 to 80) := (others => '0');
    variable r3212 : std_logic_vector(0 to 80) := (others => '0');
    variable r3210 : std_logic_vector(0 to 0) := (others => '0');
    variable r3207 : std_logic_vector(0 to 80) := (others => '0');
    variable r3203 : std_logic_vector(0 to 80) := (others => '0');
    variable r3195 : std_logic_vector(0 to 80) := (others => '0');
    variable b3191 : boolean := false;
    variable r3186 : std_logic_vector(0 to 80) := (others => '0');
    variable b3182 : boolean := false;
    variable r3177 : std_logic_vector(0 to 80) := (others => '0');
    variable b3173 : boolean := false;
    variable r3170 : std_logic_vector(0 to 1) := (others => '0');
    variable r3166 : std_logic_vector(0 to 80) := (others => '0');
    variable r3164 : std_logic_vector(0 to 7) := (others => '0');
    variable r3159 : std_logic_vector(0 to 7) := (others => '0');
    variable r3153 : std_logic_vector(0 to 7) := (others => '0');
    variable b3150 : boolean := false;
    variable r3146 : std_logic_vector(0 to 7) := (others => '0');
    variable b3143 : boolean := false;
    variable r3139 : std_logic_vector(0 to 7) := (others => '0');
    variable b3136 : boolean := false;
    variable r3134 : std_logic_vector(0 to 7) := (others => '0');
    variable r3132 : std_logic_vector(0 to 1) := (others => '0');
    variable r3128 : std_logic_vector(0 to 80) := (others => '0');
    variable r3125 : std_logic_vector(0 to 7) := (others => '0');
    variable r3119 : std_logic_vector(0 to 7) := (others => '0');
    variable b3116 : boolean := false;
    variable r3112 : std_logic_vector(0 to 7) := (others => '0');
    variable b3109 : boolean := false;
    variable r3105 : std_logic_vector(0 to 7) := (others => '0');
    variable b3102 : boolean := false;
    variable r3100 : std_logic_vector(0 to 7) := (others => '0');
    variable r3098 : std_logic_vector(0 to 1) := (others => '0');
    variable r3094 : std_logic_vector(0 to 80) := (others => '0');
    variable b3092 : boolean := false;
    variable b3090 : boolean := false;
    variable b3088 : boolean := false;
    variable b3086 : boolean := false;
    variable b3084 : boolean := false;
    variable b3082 : boolean := false;
    variable b3080 : boolean := false;
    variable b3078 : boolean := false;
    variable b3076 : boolean := false;
    variable r3074 : std_logic_vector(0 to 0) := (others => '0');
    variable r3072 : std_logic_vector(0 to 0) := (others => '0');
    variable r3070 : std_logic_vector(0 to 0) := (others => '0');
    variable r3068 : std_logic_vector(0 to 0) := (others => '0');
    variable r3066 : std_logic_vector(0 to 0) := (others => '0');
    variable r3064 : std_logic_vector(0 to 0) := (others => '0');
    variable r3062 : std_logic_vector(0 to 0) := (others => '0');
    variable r3060 : std_logic_vector(0 to 0) := (others => '0');
    variable b3058 : boolean := false;
    variable r3053 : std_logic_vector(0 to 80) := (others => '0');
    variable r3049 : std_logic_vector(0 to 80) := (others => '0');
    variable r3047 : std_logic_vector(0 to 9) := (others => '0');
    variable r3043 : std_logic_vector(0 to 17) := (others => '0');
    variable r3040 : std_logic_vector(0 to 80) := (others => '0');
    variable r3037 : std_logic_vector(0 to 80) := (others => '0');
    variable r3035 : std_logic_vector(0 to 0) := (others => '0');
    variable r3033 : std_logic_vector(0 to 7) := (others => '0');
    variable r3029 : std_logic_vector(0 to 80) := (others => '0');
    variable r3026 : std_logic_vector(0 to 80) := (others => '0');
    variable r3024 : std_logic_vector(0 to 0) := (others => '0');
    variable r3021 : std_logic_vector(0 to 80) := (others => '0');
    variable r3017 : std_logic_vector(0 to 80) := (others => '0');
    variable r3009 : std_logic_vector(0 to 80) := (others => '0');
    variable b3005 : boolean := false;
    variable r3000 : std_logic_vector(0 to 80) := (others => '0');
    variable b2996 : boolean := false;
    variable r2991 : std_logic_vector(0 to 80) := (others => '0');
    variable b2987 : boolean := false;
    variable r2984 : std_logic_vector(0 to 1) := (others => '0');
    variable r2980 : std_logic_vector(0 to 80) := (others => '0');
    variable r2978 : std_logic_vector(0 to 7) := (others => '0');
    variable r2973 : std_logic_vector(0 to 7) := (others => '0');
    variable r2967 : std_logic_vector(0 to 7) := (others => '0');
    variable b2964 : boolean := false;
    variable r2960 : std_logic_vector(0 to 7) := (others => '0');
    variable b2957 : boolean := false;
    variable r2953 : std_logic_vector(0 to 7) := (others => '0');
    variable b2950 : boolean := false;
    variable r2948 : std_logic_vector(0 to 7) := (others => '0');
    variable r2946 : std_logic_vector(0 to 1) := (others => '0');
    variable r2942 : std_logic_vector(0 to 80) := (others => '0');
    variable r2939 : std_logic_vector(0 to 7) := (others => '0');
    variable r2933 : std_logic_vector(0 to 7) := (others => '0');
    variable b2930 : boolean := false;
    variable r2926 : std_logic_vector(0 to 7) := (others => '0');
    variable b2923 : boolean := false;
    variable r2919 : std_logic_vector(0 to 7) := (others => '0');
    variable b2916 : boolean := false;
    variable r2914 : std_logic_vector(0 to 7) := (others => '0');
    variable r2912 : std_logic_vector(0 to 1) := (others => '0');
    variable r2908 : std_logic_vector(0 to 80) := (others => '0');
    variable b2906 : boolean := false;
    variable b2904 : boolean := false;
    variable b2902 : boolean := false;
    variable b2900 : boolean := false;
    variable b2898 : boolean := false;
    variable b2896 : boolean := false;
    variable b2894 : boolean := false;
    variable b2892 : boolean := false;
    variable b2890 : boolean := false;
    variable r2888 : std_logic_vector(0 to 0) := (others => '0');
    variable r2886 : std_logic_vector(0 to 0) := (others => '0');
    variable r2884 : std_logic_vector(0 to 0) := (others => '0');
    variable r2882 : std_logic_vector(0 to 0) := (others => '0');
    variable r2880 : std_logic_vector(0 to 0) := (others => '0');
    variable r2878 : std_logic_vector(0 to 0) := (others => '0');
    variable r2876 : std_logic_vector(0 to 0) := (others => '0');
    variable r2874 : std_logic_vector(0 to 0) := (others => '0');
    variable b2872 : boolean := false;
    variable r2867 : std_logic_vector(0 to 80) := (others => '0');
    variable r2863 : std_logic_vector(0 to 80) := (others => '0');
    variable r2861 : std_logic_vector(0 to 9) := (others => '0');
    variable r2857 : std_logic_vector(0 to 17) := (others => '0');
    variable r2854 : std_logic_vector(0 to 80) := (others => '0');
    variable r2851 : std_logic_vector(0 to 80) := (others => '0');
    variable r2849 : std_logic_vector(0 to 0) := (others => '0');
    variable r2847 : std_logic_vector(0 to 7) := (others => '0');
    variable r2843 : std_logic_vector(0 to 80) := (others => '0');
    variable r2840 : std_logic_vector(0 to 80) := (others => '0');
    variable r2838 : std_logic_vector(0 to 0) := (others => '0');
    variable r2835 : std_logic_vector(0 to 80) := (others => '0');
    variable r2831 : std_logic_vector(0 to 80) := (others => '0');
    variable r2823 : std_logic_vector(0 to 80) := (others => '0');
    variable b2819 : boolean := false;
    variable r2814 : std_logic_vector(0 to 80) := (others => '0');
    variable b2810 : boolean := false;
    variable r2805 : std_logic_vector(0 to 80) := (others => '0');
    variable b2801 : boolean := false;
    variable r2798 : std_logic_vector(0 to 1) := (others => '0');
    variable r2794 : std_logic_vector(0 to 80) := (others => '0');
    variable r2792 : std_logic_vector(0 to 7) := (others => '0');
    variable r2787 : std_logic_vector(0 to 7) := (others => '0');
    variable r2781 : std_logic_vector(0 to 7) := (others => '0');
    variable b2778 : boolean := false;
    variable r2774 : std_logic_vector(0 to 7) := (others => '0');
    variable b2771 : boolean := false;
    variable r2767 : std_logic_vector(0 to 7) := (others => '0');
    variable b2764 : boolean := false;
    variable r2762 : std_logic_vector(0 to 7) := (others => '0');
    variable r2760 : std_logic_vector(0 to 1) := (others => '0');
    variable r2756 : std_logic_vector(0 to 80) := (others => '0');
    variable r2753 : std_logic_vector(0 to 7) := (others => '0');
    variable r2747 : std_logic_vector(0 to 7) := (others => '0');
    variable b2744 : boolean := false;
    variable r2740 : std_logic_vector(0 to 7) := (others => '0');
    variable b2737 : boolean := false;
    variable r2733 : std_logic_vector(0 to 7) := (others => '0');
    variable b2730 : boolean := false;
    variable r2728 : std_logic_vector(0 to 7) := (others => '0');
    variable r2726 : std_logic_vector(0 to 1) := (others => '0');
    variable r2722 : std_logic_vector(0 to 80) := (others => '0');
    variable b2720 : boolean := false;
    variable b2718 : boolean := false;
    variable b2716 : boolean := false;
    variable b2714 : boolean := false;
    variable b2712 : boolean := false;
    variable b2710 : boolean := false;
    variable b2708 : boolean := false;
    variable b2706 : boolean := false;
    variable b2704 : boolean := false;
    variable r2702 : std_logic_vector(0 to 0) := (others => '0');
    variable r2700 : std_logic_vector(0 to 0) := (others => '0');
    variable r2698 : std_logic_vector(0 to 0) := (others => '0');
    variable r2696 : std_logic_vector(0 to 0) := (others => '0');
    variable r2694 : std_logic_vector(0 to 0) := (others => '0');
    variable r2692 : std_logic_vector(0 to 0) := (others => '0');
    variable r2690 : std_logic_vector(0 to 0) := (others => '0');
    variable r2688 : std_logic_vector(0 to 0) := (others => '0');
    variable b2686 : boolean := false;
    variable r2681 : std_logic_vector(0 to 80) := (others => '0');
    variable r2677 : std_logic_vector(0 to 80) := (others => '0');
    variable r2675 : std_logic_vector(0 to 9) := (others => '0');
    variable r2671 : std_logic_vector(0 to 17) := (others => '0');
    variable r2668 : std_logic_vector(0 to 80) := (others => '0');
    variable r2664 : std_logic_vector(0 to 80) := (others => '0');
    variable r2656 : std_logic_vector(0 to 80) := (others => '0');
    variable b2652 : boolean := false;
    variable r2647 : std_logic_vector(0 to 80) := (others => '0');
    variable b2643 : boolean := false;
    variable r2638 : std_logic_vector(0 to 80) := (others => '0');
    variable b2634 : boolean := false;
    variable r2631 : std_logic_vector(0 to 1) := (others => '0');
    variable r2627 : std_logic_vector(0 to 80) := (others => '0');
    variable r2624 : std_logic_vector(0 to 7) := (others => '0');
    variable r2618 : std_logic_vector(0 to 7) := (others => '0');
    variable b2615 : boolean := false;
    variable r2611 : std_logic_vector(0 to 7) := (others => '0');
    variable b2608 : boolean := false;
    variable r2604 : std_logic_vector(0 to 7) := (others => '0');
    variable b2601 : boolean := false;
    variable r2599 : std_logic_vector(0 to 7) := (others => '0');
    variable r2597 : std_logic_vector(0 to 1) := (others => '0');
    variable r2593 : std_logic_vector(0 to 80) := (others => '0');
    variable b2591 : boolean := false;
    variable b2589 : boolean := false;
    variable b2587 : boolean := false;
    variable b2585 : boolean := false;
    variable b2583 : boolean := false;
    variable b2581 : boolean := false;
    variable b2579 : boolean := false;
    variable b2577 : boolean := false;
    variable b2575 : boolean := false;
    variable r2573 : std_logic_vector(0 to 0) := (others => '0');
    variable r2571 : std_logic_vector(0 to 0) := (others => '0');
    variable r2569 : std_logic_vector(0 to 0) := (others => '0');
    variable r2567 : std_logic_vector(0 to 0) := (others => '0');
    variable r2565 : std_logic_vector(0 to 0) := (others => '0');
    variable r2563 : std_logic_vector(0 to 0) := (others => '0');
    variable r2561 : std_logic_vector(0 to 0) := (others => '0');
    variable r2559 : std_logic_vector(0 to 0) := (others => '0');
    variable b2557 : boolean := false;
    variable r2552 : std_logic_vector(0 to 80) := (others => '0');
    variable r2548 : std_logic_vector(0 to 80) := (others => '0');
    variable r2546 : std_logic_vector(0 to 9) := (others => '0');
    variable r2542 : std_logic_vector(0 to 17) := (others => '0');
    variable r2539 : std_logic_vector(0 to 80) := (others => '0');
    variable r2535 : std_logic_vector(0 to 80) := (others => '0');
    variable r2527 : std_logic_vector(0 to 80) := (others => '0');
    variable b2523 : boolean := false;
    variable r2518 : std_logic_vector(0 to 80) := (others => '0');
    variable b2514 : boolean := false;
    variable r2509 : std_logic_vector(0 to 80) := (others => '0');
    variable b2505 : boolean := false;
    variable r2502 : std_logic_vector(0 to 1) := (others => '0');
    variable r2498 : std_logic_vector(0 to 80) := (others => '0');
    variable r2495 : std_logic_vector(0 to 80) := (others => '0');
    variable r2491 : std_logic_vector(0 to 80) := (others => '0');
    variable b2486 : boolean := false;
    variable b2484 : boolean := false;
    variable r2482 : std_logic_vector(0 to 7) := (others => '0');
    variable r2480 : std_logic_vector(0 to 0) := (others => '0');
    variable r2478 : std_logic_vector(0 to 7) := (others => '0');
    variable b2472 : boolean := false;
    variable b2470 : boolean := false;
    variable r2468 : std_logic_vector(0 to 7) := (others => '0');
    variable r2466 : std_logic_vector(0 to 0) := (others => '0');
    variable r2464 : std_logic_vector(0 to 0) := (others => '0');
    variable r2461 : std_logic_vector(0 to 8) := (others => '0');
    variable r2456 : std_logic_vector(0 to 0) := (others => '0');
    variable r2453 : std_logic_vector(0 to 80) := (others => '0');
    variable r2450 : std_logic_vector(0 to 7) := (others => '0');
    variable r2444 : std_logic_vector(0 to 7) := (others => '0');
    variable b2441 : boolean := false;
    variable r2437 : std_logic_vector(0 to 7) := (others => '0');
    variable b2434 : boolean := false;
    variable r2430 : std_logic_vector(0 to 7) := (others => '0');
    variable b2427 : boolean := false;
    variable r2425 : std_logic_vector(0 to 7) := (others => '0');
    variable r2423 : std_logic_vector(0 to 1) := (others => '0');
    variable r2419 : std_logic_vector(0 to 80) := (others => '0');
    variable r2416 : std_logic_vector(0 to 7) := (others => '0');
    variable r2410 : std_logic_vector(0 to 7) := (others => '0');
    variable b2407 : boolean := false;
    variable r2403 : std_logic_vector(0 to 7) := (others => '0');
    variable b2400 : boolean := false;
    variable r2396 : std_logic_vector(0 to 7) := (others => '0');
    variable b2393 : boolean := false;
    variable r2391 : std_logic_vector(0 to 7) := (others => '0');
    variable r2389 : std_logic_vector(0 to 1) := (others => '0');
    variable r2385 : std_logic_vector(0 to 80) := (others => '0');
    variable b2383 : boolean := false;
    variable b2381 : boolean := false;
    variable b2379 : boolean := false;
    variable b2377 : boolean := false;
    variable b2375 : boolean := false;
    variable b2373 : boolean := false;
    variable b2371 : boolean := false;
    variable b2369 : boolean := false;
    variable b2367 : boolean := false;
    variable r2365 : std_logic_vector(0 to 0) := (others => '0');
    variable r2363 : std_logic_vector(0 to 0) := (others => '0');
    variable r2361 : std_logic_vector(0 to 0) := (others => '0');
    variable r2359 : std_logic_vector(0 to 0) := (others => '0');
    variable r2357 : std_logic_vector(0 to 0) := (others => '0');
    variable r2355 : std_logic_vector(0 to 0) := (others => '0');
    variable r2353 : std_logic_vector(0 to 0) := (others => '0');
    variable r2351 : std_logic_vector(0 to 0) := (others => '0');
    variable b2349 : boolean := false;
    variable r2344 : std_logic_vector(0 to 80) := (others => '0');
    variable r2340 : std_logic_vector(0 to 80) := (others => '0');
    variable r2338 : std_logic_vector(0 to 9) := (others => '0');
    variable r2334 : std_logic_vector(0 to 17) := (others => '0');
    variable r2331 : std_logic_vector(0 to 80) := (others => '0');
    variable r2327 : std_logic_vector(0 to 80) := (others => '0');
    variable r2319 : std_logic_vector(0 to 80) := (others => '0');
    variable b2315 : boolean := false;
    variable r2310 : std_logic_vector(0 to 80) := (others => '0');
    variable b2306 : boolean := false;
    variable r2301 : std_logic_vector(0 to 80) := (others => '0');
    variable b2297 : boolean := false;
    variable r2294 : std_logic_vector(0 to 1) := (others => '0');
    variable r2290 : std_logic_vector(0 to 80) := (others => '0');
    variable r2287 : std_logic_vector(0 to 80) := (others => '0');
    variable r2283 : std_logic_vector(0 to 80) := (others => '0');
    variable b2278 : boolean := false;
    variable b2276 : boolean := false;
    variable r2274 : std_logic_vector(0 to 7) := (others => '0');
    variable r2272 : std_logic_vector(0 to 0) := (others => '0');
    variable r2270 : std_logic_vector(0 to 7) := (others => '0');
    variable b2264 : boolean := false;
    variable b2262 : boolean := false;
    variable r2260 : std_logic_vector(0 to 7) := (others => '0');
    variable r2258 : std_logic_vector(0 to 0) := (others => '0');
    variable r2256 : std_logic_vector(0 to 0) := (others => '0');
    variable r2253 : std_logic_vector(0 to 8) := (others => '0');
    variable r2251 : std_logic_vector(0 to 0) := (others => '0');
    variable r2246 : std_logic_vector(0 to 7) := (others => '0');
    variable r2240 : std_logic_vector(0 to 7) := (others => '0');
    variable b2237 : boolean := false;
    variable r2233 : std_logic_vector(0 to 7) := (others => '0');
    variable b2230 : boolean := false;
    variable r2226 : std_logic_vector(0 to 7) := (others => '0');
    variable b2223 : boolean := false;
    variable r2221 : std_logic_vector(0 to 7) := (others => '0');
    variable r2219 : std_logic_vector(0 to 1) := (others => '0');
    variable r2215 : std_logic_vector(0 to 80) := (others => '0');
    variable r2212 : std_logic_vector(0 to 7) := (others => '0');
    variable r2206 : std_logic_vector(0 to 7) := (others => '0');
    variable b2203 : boolean := false;
    variable r2199 : std_logic_vector(0 to 7) := (others => '0');
    variable b2196 : boolean := false;
    variable r2192 : std_logic_vector(0 to 7) := (others => '0');
    variable b2189 : boolean := false;
    variable r2187 : std_logic_vector(0 to 7) := (others => '0');
    variable r2185 : std_logic_vector(0 to 1) := (others => '0');
    variable r2181 : std_logic_vector(0 to 80) := (others => '0');
    variable b2179 : boolean := false;
    variable b2177 : boolean := false;
    variable b2175 : boolean := false;
    variable b2173 : boolean := false;
    variable b2171 : boolean := false;
    variable b2169 : boolean := false;
    variable b2167 : boolean := false;
    variable b2165 : boolean := false;
    variable b2163 : boolean := false;
    variable r2161 : std_logic_vector(0 to 0) := (others => '0');
    variable r2159 : std_logic_vector(0 to 0) := (others => '0');
    variable r2157 : std_logic_vector(0 to 0) := (others => '0');
    variable r2155 : std_logic_vector(0 to 0) := (others => '0');
    variable r2153 : std_logic_vector(0 to 0) := (others => '0');
    variable r2151 : std_logic_vector(0 to 0) := (others => '0');
    variable r2149 : std_logic_vector(0 to 0) := (others => '0');
    variable r2147 : std_logic_vector(0 to 0) := (others => '0');
    variable b2145 : boolean := false;
    variable r2140 : std_logic_vector(0 to 80) := (others => '0');
    variable r2136 : std_logic_vector(0 to 80) := (others => '0');
    variable r2134 : std_logic_vector(0 to 9) := (others => '0');
    variable r2130 : std_logic_vector(0 to 17) := (others => '0');
    variable r2127 : std_logic_vector(0 to 80) := (others => '0');
    variable r2123 : std_logic_vector(0 to 80) := (others => '0');
    variable r2115 : std_logic_vector(0 to 80) := (others => '0');
    variable b2111 : boolean := false;
    variable r2106 : std_logic_vector(0 to 80) := (others => '0');
    variable b2102 : boolean := false;
    variable r2097 : std_logic_vector(0 to 80) := (others => '0');
    variable b2093 : boolean := false;
    variable r2090 : std_logic_vector(0 to 1) := (others => '0');
    variable r2086 : std_logic_vector(0 to 80) := (others => '0');
    variable r2083 : std_logic_vector(0 to 80) := (others => '0');
    variable r2079 : std_logic_vector(0 to 80) := (others => '0');
    variable b2074 : boolean := false;
    variable b2072 : boolean := false;
    variable r2070 : std_logic_vector(0 to 7) := (others => '0');
    variable r2068 : std_logic_vector(0 to 0) := (others => '0');
    variable r2066 : std_logic_vector(0 to 7) := (others => '0');
    variable b2060 : boolean := false;
    variable b2058 : boolean := false;
    variable r2056 : std_logic_vector(0 to 7) := (others => '0');
    variable r2054 : std_logic_vector(0 to 0) := (others => '0');
    variable r2052 : std_logic_vector(0 to 0) := (others => '0');
    variable r2049 : std_logic_vector(0 to 8) := (others => '0');
    variable r2044 : std_logic_vector(0 to 0) := (others => '0');
    variable r2041 : std_logic_vector(0 to 80) := (others => '0');
    variable r2038 : std_logic_vector(0 to 7) := (others => '0');
    variable r2032 : std_logic_vector(0 to 7) := (others => '0');
    variable b2029 : boolean := false;
    variable r2025 : std_logic_vector(0 to 7) := (others => '0');
    variable b2022 : boolean := false;
    variable r2018 : std_logic_vector(0 to 7) := (others => '0');
    variable b2015 : boolean := false;
    variable r2013 : std_logic_vector(0 to 7) := (others => '0');
    variable r2011 : std_logic_vector(0 to 1) := (others => '0');
    variable r2007 : std_logic_vector(0 to 80) := (others => '0');
    variable r2004 : std_logic_vector(0 to 7) := (others => '0');
    variable r1998 : std_logic_vector(0 to 7) := (others => '0');
    variable b1995 : boolean := false;
    variable r1991 : std_logic_vector(0 to 7) := (others => '0');
    variable b1988 : boolean := false;
    variable r1984 : std_logic_vector(0 to 7) := (others => '0');
    variable b1981 : boolean := false;
    variable r1979 : std_logic_vector(0 to 7) := (others => '0');
    variable r1977 : std_logic_vector(0 to 1) := (others => '0');
    variable r1973 : std_logic_vector(0 to 80) := (others => '0');
    variable b1971 : boolean := false;
    variable b1969 : boolean := false;
    variable b1967 : boolean := false;
    variable b1965 : boolean := false;
    variable b1963 : boolean := false;
    variable b1961 : boolean := false;
    variable b1959 : boolean := false;
    variable b1957 : boolean := false;
    variable b1955 : boolean := false;
    variable r1953 : std_logic_vector(0 to 0) := (others => '0');
    variable r1951 : std_logic_vector(0 to 0) := (others => '0');
    variable r1949 : std_logic_vector(0 to 0) := (others => '0');
    variable r1947 : std_logic_vector(0 to 0) := (others => '0');
    variable r1945 : std_logic_vector(0 to 0) := (others => '0');
    variable r1943 : std_logic_vector(0 to 0) := (others => '0');
    variable r1941 : std_logic_vector(0 to 0) := (others => '0');
    variable r1939 : std_logic_vector(0 to 0) := (others => '0');
    variable b1937 : boolean := false;
    variable r1932 : std_logic_vector(0 to 80) := (others => '0');
    variable r1928 : std_logic_vector(0 to 80) := (others => '0');
    variable r1926 : std_logic_vector(0 to 9) := (others => '0');
    variable r1922 : std_logic_vector(0 to 17) := (others => '0');
    variable r1919 : std_logic_vector(0 to 80) := (others => '0');
    variable r1915 : std_logic_vector(0 to 80) := (others => '0');
    variable r1907 : std_logic_vector(0 to 80) := (others => '0');
    variable b1903 : boolean := false;
    variable r1898 : std_logic_vector(0 to 80) := (others => '0');
    variable b1894 : boolean := false;
    variable r1889 : std_logic_vector(0 to 80) := (others => '0');
    variable b1885 : boolean := false;
    variable r1882 : std_logic_vector(0 to 1) := (others => '0');
    variable r1878 : std_logic_vector(0 to 80) := (others => '0');
    variable r1875 : std_logic_vector(0 to 80) := (others => '0');
    variable r1871 : std_logic_vector(0 to 80) := (others => '0');
    variable b1866 : boolean := false;
    variable b1864 : boolean := false;
    variable r1862 : std_logic_vector(0 to 7) := (others => '0');
    variable r1860 : std_logic_vector(0 to 0) := (others => '0');
    variable r1858 : std_logic_vector(0 to 7) := (others => '0');
    variable b1852 : boolean := false;
    variable b1850 : boolean := false;
    variable r1848 : std_logic_vector(0 to 7) := (others => '0');
    variable r1846 : std_logic_vector(0 to 0) := (others => '0');
    variable r1844 : std_logic_vector(0 to 0) := (others => '0');
    variable r1841 : std_logic_vector(0 to 8) := (others => '0');
    variable r1839 : std_logic_vector(0 to 0) := (others => '0');
    variable r1834 : std_logic_vector(0 to 7) := (others => '0');
    variable r1828 : std_logic_vector(0 to 7) := (others => '0');
    variable b1825 : boolean := false;
    variable r1821 : std_logic_vector(0 to 7) := (others => '0');
    variable b1818 : boolean := false;
    variable r1814 : std_logic_vector(0 to 7) := (others => '0');
    variable b1811 : boolean := false;
    variable r1809 : std_logic_vector(0 to 7) := (others => '0');
    variable r1807 : std_logic_vector(0 to 1) := (others => '0');
    variable r1803 : std_logic_vector(0 to 80) := (others => '0');
    variable r1800 : std_logic_vector(0 to 7) := (others => '0');
    variable r1794 : std_logic_vector(0 to 7) := (others => '0');
    variable b1791 : boolean := false;
    variable r1787 : std_logic_vector(0 to 7) := (others => '0');
    variable b1784 : boolean := false;
    variable r1780 : std_logic_vector(0 to 7) := (others => '0');
    variable b1777 : boolean := false;
    variable r1775 : std_logic_vector(0 to 7) := (others => '0');
    variable r1773 : std_logic_vector(0 to 1) := (others => '0');
    variable r1769 : std_logic_vector(0 to 80) := (others => '0');
    variable b1767 : boolean := false;
    variable b1765 : boolean := false;
    variable b1763 : boolean := false;
    variable b1761 : boolean := false;
    variable b1759 : boolean := false;
    variable b1757 : boolean := false;
    variable b1755 : boolean := false;
    variable b1753 : boolean := false;
    variable b1751 : boolean := false;
    variable r1749 : std_logic_vector(0 to 0) := (others => '0');
    variable r1747 : std_logic_vector(0 to 0) := (others => '0');
    variable r1745 : std_logic_vector(0 to 0) := (others => '0');
    variable r1743 : std_logic_vector(0 to 0) := (others => '0');
    variable r1741 : std_logic_vector(0 to 0) := (others => '0');
    variable r1739 : std_logic_vector(0 to 0) := (others => '0');
    variable r1737 : std_logic_vector(0 to 0) := (others => '0');
    variable r1735 : std_logic_vector(0 to 0) := (others => '0');
    variable b1733 : boolean := false;
    variable r1728 : std_logic_vector(0 to 80) := (others => '0');
    variable r1724 : std_logic_vector(0 to 80) := (others => '0');
    variable r1722 : std_logic_vector(0 to 9) := (others => '0');
    variable r1718 : std_logic_vector(0 to 17) := (others => '0');
    variable r1715 : std_logic_vector(0 to 80) := (others => '0');
    variable r1712 : std_logic_vector(0 to 80) := (others => '0');
    variable r1710 : std_logic_vector(0 to 17) := (others => '0');
    variable r1705 : std_logic_vector(0 to 80) := (others => '0');
    variable r1703 : std_logic_vector(0 to 17) := (others => '0');
    variable r1700 : std_logic_vector(0 to 80) := (others => '0');
    variable r1697 : std_logic_vector(0 to 80) := (others => '0');
    variable r1695 : std_logic_vector(0 to 17) := (others => '0');
    variable r1690 : std_logic_vector(0 to 80) := (others => '0');
    variable r1688 : std_logic_vector(0 to 17) := (others => '0');
    variable r1685 : std_logic_vector(0 to 80) := (others => '0');
    variable r1682 : std_logic_vector(0 to 80) := (others => '0');
    variable r1680 : std_logic_vector(0 to 17) := (others => '0');
    variable r1678 : std_logic_vector(0 to 0) := (others => '0');
    variable r1674 : std_logic_vector(0 to 80) := (others => '0');
    variable r1672 : std_logic_vector(0 to 17) := (others => '0');
    variable r1669 : std_logic_vector(0 to 80) := (others => '0');
    variable r1666 : std_logic_vector(0 to 7) := (others => '0');
    variable r1660 : std_logic_vector(0 to 7) := (others => '0');
    variable b1657 : boolean := false;
    variable r1653 : std_logic_vector(0 to 7) := (others => '0');
    variable b1650 : boolean := false;
    variable r1646 : std_logic_vector(0 to 7) := (others => '0');
    variable b1643 : boolean := false;
    variable r1641 : std_logic_vector(0 to 7) := (others => '0');
    variable r1639 : std_logic_vector(0 to 1) := (others => '0');
    variable r1635 : std_logic_vector(0 to 80) := (others => '0');
    variable r1632 : std_logic_vector(0 to 7) := (others => '0');
    variable r1626 : std_logic_vector(0 to 7) := (others => '0');
    variable b1623 : boolean := false;
    variable r1619 : std_logic_vector(0 to 7) := (others => '0');
    variable b1616 : boolean := false;
    variable r1612 : std_logic_vector(0 to 7) := (others => '0');
    variable b1609 : boolean := false;
    variable r1607 : std_logic_vector(0 to 7) := (others => '0');
    variable r1605 : std_logic_vector(0 to 1) := (others => '0');
    variable r1601 : std_logic_vector(0 to 80) := (others => '0');
    variable b1599 : boolean := false;
    variable b1597 : boolean := false;
    variable b1595 : boolean := false;
    variable b1593 : boolean := false;
    variable b1591 : boolean := false;
    variable b1589 : boolean := false;
    variable b1587 : boolean := false;
    variable b1585 : boolean := false;
    variable b1583 : boolean := false;
    variable r1581 : std_logic_vector(0 to 0) := (others => '0');
    variable r1579 : std_logic_vector(0 to 0) := (others => '0');
    variable r1577 : std_logic_vector(0 to 0) := (others => '0');
    variable r1575 : std_logic_vector(0 to 0) := (others => '0');
    variable r1573 : std_logic_vector(0 to 0) := (others => '0');
    variable r1571 : std_logic_vector(0 to 0) := (others => '0');
    variable r1569 : std_logic_vector(0 to 0) := (others => '0');
    variable r1567 : std_logic_vector(0 to 0) := (others => '0');
    variable b1565 : boolean := false;
    variable r1559 : std_logic_vector(0 to 80) := (others => '0');
    variable r1551 : std_logic_vector(0 to 80) := (others => '0');
    variable b1547 : boolean := false;
    variable r1542 : std_logic_vector(0 to 80) := (others => '0');
    variable b1538 : boolean := false;
    variable r1533 : std_logic_vector(0 to 80) := (others => '0');
    variable b1529 : boolean := false;
    variable r1526 : std_logic_vector(0 to 1) := (others => '0');
    variable r1522 : std_logic_vector(0 to 80) := (others => '0');
    variable r1520 : std_logic_vector(0 to 7) := (others => '0');
    variable r1517 : std_logic_vector(0 to 9) := (others => '0');
    variable r1514 : std_logic_vector(0 to 80) := (others => '0');
    variable r1511 : std_logic_vector(0 to 80) := (others => '0');
    variable r1507 : std_logic_vector(0 to 80) := (others => '0');
    variable r1505 : std_logic_vector(0 to 9) := (others => '0');
    variable r1501 : std_logic_vector(0 to 17) := (others => '0');
    variable r1498 : std_logic_vector(0 to 80) := (others => '0');
    variable r1495 : std_logic_vector(0 to 80) := (others => '0');
    variable r1493 : std_logic_vector(0 to 17) := (others => '0');
    variable r1488 : std_logic_vector(0 to 80) := (others => '0');
    variable r1486 : std_logic_vector(0 to 17) := (others => '0');
    variable r1483 : std_logic_vector(0 to 80) := (others => '0');
    variable r1480 : std_logic_vector(0 to 80) := (others => '0');
    variable r1478 : std_logic_vector(0 to 17) := (others => '0');
    variable r1476 : std_logic_vector(0 to 0) := (others => '0');
    variable r1472 : std_logic_vector(0 to 80) := (others => '0');
    variable r1470 : std_logic_vector(0 to 17) := (others => '0');
    variable r1467 : std_logic_vector(0 to 80) := (others => '0');
    variable r1464 : std_logic_vector(0 to 7) := (others => '0');
    variable r1458 : std_logic_vector(0 to 7) := (others => '0');
    variable b1455 : boolean := false;
    variable r1451 : std_logic_vector(0 to 7) := (others => '0');
    variable b1448 : boolean := false;
    variable r1444 : std_logic_vector(0 to 7) := (others => '0');
    variable b1441 : boolean := false;
    variable r1439 : std_logic_vector(0 to 7) := (others => '0');
    variable r1437 : std_logic_vector(0 to 1) := (others => '0');
    variable r1433 : std_logic_vector(0 to 80) := (others => '0');
    variable b1431 : boolean := false;
    variable b1429 : boolean := false;
    variable b1427 : boolean := false;
    variable b1425 : boolean := false;
    variable b1423 : boolean := false;
    variable b1421 : boolean := false;
    variable b1419 : boolean := false;
    variable b1417 : boolean := false;
    variable b1415 : boolean := false;
    variable r1413 : std_logic_vector(0 to 0) := (others => '0');
    variable r1411 : std_logic_vector(0 to 0) := (others => '0');
    variable r1409 : std_logic_vector(0 to 0) := (others => '0');
    variable r1407 : std_logic_vector(0 to 0) := (others => '0');
    variable r1405 : std_logic_vector(0 to 0) := (others => '0');
    variable r1403 : std_logic_vector(0 to 0) := (others => '0');
    variable r1401 : std_logic_vector(0 to 0) := (others => '0');
    variable r1399 : std_logic_vector(0 to 0) := (others => '0');
    variable b1397 : boolean := false;
    variable r1386 : std_logic_vector(0 to 80) := (others => '0');
    variable r1352 : std_logic_vector(0 to 80) := (others => '0');
    variable r1351 : std_logic_vector(0 to 7) := (others => '0');
    variable r1350 : std_logic_vector(0 to 80) := (others => '0');
    variable r1343 : std_logic_vector(0 to 80) := (others => '0');
    variable r1309 : std_logic_vector(0 to 80) := (others => '0');
    variable r1308 : std_logic_vector(0 to 7) := (others => '0');
    variable r1307 : std_logic_vector(0 to 80) := (others => '0');
    variable b1304 : boolean := false;
    variable r1299 : std_logic_vector(0 to 80) := (others => '0');
    variable r1265 : std_logic_vector(0 to 80) := (others => '0');
    variable r1264 : std_logic_vector(0 to 7) := (others => '0');
    variable r1263 : std_logic_vector(0 to 80) := (others => '0');
    variable b1260 : boolean := false;
    variable r1255 : std_logic_vector(0 to 80) := (others => '0');
    variable r1221 : std_logic_vector(0 to 80) := (others => '0');
    variable r1220 : std_logic_vector(0 to 7) := (others => '0');
    variable r1219 : std_logic_vector(0 to 80) := (others => '0');
    variable b1216 : boolean := false;
    variable r1213 : std_logic_vector(0 to 1) := (others => '0');
    variable r1209 : std_logic_vector(0 to 80) := (others => '0');
    variable r1207 : std_logic_vector(0 to 7) := (others => '0');
    variable r1204 : std_logic_vector(0 to 9) := (others => '0');
    variable r1201 : std_logic_vector(0 to 80) := (others => '0');
    variable b1199 : boolean := false;
    variable r1194 : std_logic_vector(0 to 80) := (others => '0');
    variable r1190 : std_logic_vector(0 to 80) := (others => '0');
    variable r1188 : std_logic_vector(0 to 9) := (others => '0');
    variable r1184 : std_logic_vector(0 to 17) := (others => '0');
    variable r1181 : std_logic_vector(0 to 80) := (others => '0');
    variable r1178 : std_logic_vector(0 to 80) := (others => '0');
    variable b1173 : boolean := false;
    variable b1171 : boolean := false;
    variable r1169 : std_logic_vector(0 to 7) := (others => '0');
    variable r1167 : std_logic_vector(0 to 0) := (others => '0');
    variable r1165 : std_logic_vector(0 to 7) := (others => '0');
    variable r1163 : std_logic_vector(0 to 8) := (others => '0');
    variable r1161 : std_logic_vector(0 to 7) := (others => '0');
    variable r1127 : std_logic_vector(0 to 80) := (others => '0');
    variable r1126 : std_logic_vector(0 to 7) := (others => '0');
    variable r1125 : std_logic_vector(0 to 80) := (others => '0');
    variable r1122 : std_logic_vector(0 to 80) := (others => '0');
    variable r1119 : std_logic_vector(0 to 80) := (others => '0');
    variable r1111 : std_logic_vector(0 to 80) := (others => '0');
    variable r1109 : std_logic_vector(0 to 17) := (others => '0');
    variable r1093 : std_logic_vector(0 to 17) := (others => '0');
    variable r1092 : std_logic_vector(0 to 7) := (others => '0');
    variable r1091 : std_logic_vector(0 to 17) := (others => '0');
    variable r1087 : std_logic_vector(0 to 80) := (others => '0');
    variable r1085 : std_logic_vector(0 to 17) := (others => '0');
    variable r1082 : std_logic_vector(0 to 80) := (others => '0');
    variable r1079 : std_logic_vector(0 to 7) := (others => '0');
    variable r1048 : std_logic_vector(0 to 7) := (others => '0');
    variable r1047 : std_logic_vector(0 to 80) := (others => '0');
    variable r1041 : std_logic_vector(0 to 7) := (others => '0');
    variable r1010 : std_logic_vector(0 to 7) := (others => '0');
    variable r1009 : std_logic_vector(0 to 80) := (others => '0');
    variable b1006 : boolean := false;
    variable r1002 : std_logic_vector(0 to 7) := (others => '0');
    variable r971 : std_logic_vector(0 to 7) := (others => '0');
    variable r970 : std_logic_vector(0 to 80) := (others => '0');
    variable b967 : boolean := false;
    variable r963 : std_logic_vector(0 to 7) := (others => '0');
    variable r932 : std_logic_vector(0 to 7) := (others => '0');
    variable r931 : std_logic_vector(0 to 80) := (others => '0');
    variable b928 : boolean := false;
    variable r926 : std_logic_vector(0 to 7) := (others => '0');
    variable r924 : std_logic_vector(0 to 1) := (others => '0');
    variable r886 : std_logic_vector(0 to 1) := (others => '0');
    variable r885 : std_logic_vector(0 to 0) := (others => '0');
    variable r884 : std_logic_vector(0 to 0) := (others => '0');
    variable r881 : std_logic_vector(0 to 80) := (others => '0');
    variable b879 : boolean := false;
    variable r874 : std_logic_vector(0 to 80) := (others => '0');
    variable r872 : std_logic_vector(0 to 17) := (others => '0');
    variable r856 : std_logic_vector(0 to 17) := (others => '0');
    variable r855 : std_logic_vector(0 to 0) := (others => '0');
    variable r854 : std_logic_vector(0 to 17) := (others => '0');
    variable r850 : std_logic_vector(0 to 80) := (others => '0');
    variable r848 : std_logic_vector(0 to 17) := (others => '0');
    variable r845 : std_logic_vector(0 to 80) := (others => '0');
    variable r842 : std_logic_vector(0 to 80) := (others => '0');
    variable r840 : std_logic_vector(0 to 17) := (others => '0');
    variable r835 : std_logic_vector(0 to 80) := (others => '0');
    variable r833 : std_logic_vector(0 to 17) := (others => '0');
    variable r830 : std_logic_vector(0 to 80) := (others => '0');
    variable r828 : std_logic_vector(0 to 7) := (others => '0');
    variable r825 : std_logic_vector(0 to 9) := (others => '0');
    variable r822 : std_logic_vector(0 to 80) := (others => '0');
    variable r819 : std_logic_vector(0 to 80) := (others => '0');
    variable r815 : std_logic_vector(0 to 80) := (others => '0');
    variable r813 : std_logic_vector(0 to 9) := (others => '0');
    variable r809 : std_logic_vector(0 to 17) := (others => '0');
    variable r806 : std_logic_vector(0 to 80) := (others => '0');
    variable r803 : std_logic_vector(0 to 80) := (others => '0');
    variable r801 : std_logic_vector(0 to 17) := (others => '0');
    variable r785 : std_logic_vector(0 to 17) := (others => '0');
    variable r784 : std_logic_vector(0 to 7) := (others => '0');
    variable r783 : std_logic_vector(0 to 17) := (others => '0');
    variable r779 : std_logic_vector(0 to 80) := (others => '0');
    variable r777 : std_logic_vector(0 to 17) := (others => '0');
    variable r774 : std_logic_vector(0 to 80) := (others => '0');
    variable r772 : std_logic_vector(0 to 7) := (others => '0');
    variable r769 : std_logic_vector(0 to 80) := (others => '0');
    variable b767 : boolean := false;
    variable b765 : boolean := false;
    variable b763 : boolean := false;
    variable b761 : boolean := false;
    variable b759 : boolean := false;
    variable b757 : boolean := false;
    variable b755 : boolean := false;
    variable b753 : boolean := false;
    variable b751 : boolean := false;
    variable r749 : std_logic_vector(0 to 0) := (others => '0');
    variable r747 : std_logic_vector(0 to 0) := (others => '0');
    variable r745 : std_logic_vector(0 to 0) := (others => '0');
    variable r743 : std_logic_vector(0 to 0) := (others => '0');
    variable r741 : std_logic_vector(0 to 0) := (others => '0');
    variable r739 : std_logic_vector(0 to 0) := (others => '0');
    variable r737 : std_logic_vector(0 to 0) := (others => '0');
    variable r735 : std_logic_vector(0 to 0) := (others => '0');
    variable b733 : boolean := false;
    variable r730 : std_logic_vector(0 to 7) := (others => '0');
    variable r719 : std_logic_vector(0 to 7) := (others => '0');
    variable r718 : std_logic_vector(0 to 9) := (others => '0');
    variable b715 : boolean := false;
    variable r710 : std_logic_vector(0 to 80) := (others => '0');
    variable r706 : std_logic_vector(0 to 80) := (others => '0');
    variable r704 : std_logic_vector(0 to 9) := (others => '0');
    variable r700 : std_logic_vector(0 to 17) := (others => '0');
    variable r697 : std_logic_vector(0 to 80) := (others => '0');
    variable r694 : std_logic_vector(0 to 80) := (others => '0');
    variable r660 : std_logic_vector(0 to 80) := (others => '0');
    variable r659 : std_logic_vector(0 to 0) := (others => '0');
    variable r658 : std_logic_vector(0 to 80) := (others => '0');
    variable r655 : std_logic_vector(0 to 80) := (others => '0');
    variable r652 : std_logic_vector(0 to 80) := (others => '0');
    variable r618 : std_logic_vector(0 to 80) := (others => '0');
    variable r617 : std_logic_vector(0 to 0) := (others => '0');
    variable r616 : std_logic_vector(0 to 80) := (others => '0');
    variable r613 : std_logic_vector(0 to 80) := (others => '0');
    variable r610 : std_logic_vector(0 to 80) := (others => '0');
    variable r576 : std_logic_vector(0 to 80) := (others => '0');
    variable r575 : std_logic_vector(0 to 7) := (others => '0');
    variable r574 : std_logic_vector(0 to 80) := (others => '0');
    variable r571 : std_logic_vector(0 to 80) := (others => '0');
    variable r569 : std_logic_vector(0 to 0) := (others => '0');
    variable r538 : std_logic_vector(0 to 0) := (others => '0');
    variable r537 : std_logic_vector(0 to 80) := (others => '0');
    variable r534 : std_logic_vector(0 to 80) := (others => '0');
    variable r532 : std_logic_vector(0 to 0) := (others => '0');
    variable r501 : std_logic_vector(0 to 0) := (others => '0');
    variable r500 : std_logic_vector(0 to 80) := (others => '0');
    variable r497 : std_logic_vector(0 to 80) := (others => '0');
    variable r495 : std_logic_vector(0 to 7) := (others => '0');
    variable r464 : std_logic_vector(0 to 7) := (others => '0');
    variable r463 : std_logic_vector(0 to 80) := (others => '0');
    variable r460 : std_logic_vector(0 to 80) := (others => '0');
    variable r457 : std_logic_vector(0 to 80) := (others => '0');
    variable r455 : std_logic_vector(0 to 0) := (others => '0');
    variable r422 : std_logic_vector(0 to 80) := (others => '0');
    variable r421 : std_logic_vector(0 to 0) := (others => '0');
    variable r420 : std_logic_vector(0 to 80) := (others => '0');
    variable r417 : std_logic_vector(0 to 80) := (others => '0');
    variable b415 : boolean := false;
    variable b413 : boolean := false;
    variable b411 : boolean := false;
    variable r409 : std_logic_vector(0 to 0) := (others => '0');
    variable r407 : std_logic_vector(0 to 0) := (others => '0');
    variable b405 : boolean := false;
    variable r402 : std_logic_vector(0 to 1) := (others => '0');
    variable r400 : std_logic_vector(0 to 0) := (others => '0');
    variable r389 : std_logic_vector(0 to 0) := (others => '0');
    variable r388 : std_logic_vector(0 to 9) := (others => '0');
    variable b380 : boolean := false;
    variable b378 : boolean := false;
    variable b376 : boolean := false;
    variable b374 : boolean := false;
    variable b372 : boolean := false;
    variable b370 : boolean := false;
    variable b368 : boolean := false;
    variable b366 : boolean := false;
    variable b364 : boolean := false;
    variable b362 : boolean := false;
    variable b360 : boolean := false;
    variable b358 : boolean := false;
    variable b356 : boolean := false;
    variable r354 : std_logic_vector(0 to 7) := (others => '0');
    variable r352 : std_logic_vector(0 to 7) := (others => '0');
    variable r350 : std_logic_vector(0 to 7) := (others => '0');
    variable r348 : std_logic_vector(0 to 7) := (others => '0');
    variable r346 : std_logic_vector(0 to 7) := (others => '0');
    variable r344 : std_logic_vector(0 to 0) := (others => '0');
    variable r342 : std_logic_vector(0 to 0) := (others => '0');
    variable r340 : std_logic_vector(0 to 7) := (others => '0');
    variable r338 : std_logic_vector(0 to 0) := (others => '0');
    variable r336 : std_logic_vector(0 to 0) := (others => '0');
    variable r334 : std_logic_vector(0 to 0) := (others => '0');
    variable r332 : std_logic_vector(0 to 17) := (others => '0');
    variable r330 : std_logic_vector(0 to 9) := (others => '0');
    variable r328 : std_logic_vector(0 to 0) := (others => '0');
    variable r325 : std_logic_vector(0 to 80) := (others => '0');
    variable r319 : std_logic_vector(0 to 80) := (others => '0');
    variable r315 : std_logic_vector(0 to 80) := (others => '0');
    variable r313 : std_logic_vector(0 to 9) := (others => '0');
    variable r309 : std_logic_vector(0 to 17) := (others => '0');
    variable r306 : std_logic_vector(0 to 80) := (others => '0');
    variable r303 : std_logic_vector(0 to 80) := (others => '0');
    variable r301 : std_logic_vector(0 to 17) := (others => '0');
    variable r298 : std_logic_vector(0 to 80) := (others => '0');
    variable r295 : std_logic_vector(0 to 80) := (others => '0');
    variable r293 : std_logic_vector(0 to 0) := (others => '0');
    variable r290 : std_logic_vector(0 to 80) := (others => '0');
    variable r287 : std_logic_vector(0 to 80) := (others => '0');
    variable r285 : std_logic_vector(0 to 0) := (others => '0');
    variable r282 : std_logic_vector(0 to 80) := (others => '0');
    variable b280 : boolean := false;
    variable r277 : std_logic_vector(0 to 0) := (others => '0');
    variable r266 : std_logic_vector(0 to 0) := (others => '0');
    variable r265 : std_logic_vector(0 to 9) := (others => '0');
    variable r262 : std_logic_vector(0 to 9) := (others => '0');
    variable r231 : std_logic_vector(0 to 9) := (others => '0');
    variable r230 : std_logic_vector(0 to 80) := (others => '0');
    variable r227 : std_logic_vector(0 to 80) := (others => '0');
    variable r222 : std_logic_vector(0 to 80) := (others => '0');
    variable r188 : std_logic_vector(0 to 80) := (others => '0');
    variable r187 : std_logic_vector(0 to 9) := (others => '0');
    variable r186 : std_logic_vector(0 to 80) := (others => '0');
    variable r183 : std_logic_vector(0 to 80) := (others => '0');
    variable r181 : std_logic_vector(0 to 9) := (others => '0');
    variable r177 : std_logic_vector(0 to 17) := (others => '0');
    variable r146 : std_logic_vector(0 to 17) := (others => '0');
    variable r145 : std_logic_vector(0 to 80) := (others => '0');
    variable r142 : std_logic_vector(0 to 80) := (others => '0');
    variable r139 : std_logic_vector(0 to 80) := (others => '0');
    variable r137 : std_logic_vector(0 to 17) := (others => '0');
    variable r128 : std_logic_vector(0 to 17) := (others => '0');
    variable r94 : std_logic_vector(0 to 80) := (others => '0');
    variable r93 : std_logic_vector(0 to 17) := (others => '0');
    variable r92 : std_logic_vector(0 to 80) := (others => '0');
    variable r89 : std_logic_vector(0 to 80) := (others => '0');
    variable r86 : std_logic_vector(0 to 80) := (others => '0');
    variable r84 : std_logic_vector(0 to 0) := (others => '0');
    variable r51 : std_logic_vector(0 to 80) := (others => '0');
    variable r50 : std_logic_vector(0 to 0) := (others => '0');
    variable r49 : std_logic_vector(0 to 80) := (others => '0');
    variable r46 : std_logic_vector(0 to 80) := (others => '0');
    variable r43 : std_logic_vector(0 to 80) := (others => '0');
    variable r41 : std_logic_vector(0 to 0) := (others => '0');
    variable r8 : std_logic_vector(0 to 80) := (others => '0');
    variable r7 : std_logic_vector(0 to 0) := (others => '0');
    variable r6 : std_logic_vector(0 to 80) := (others => '0');
    variable r3 : std_logic_vector(0 to 80) := (others => '0');
    variable EMPTY : std_logic_vector(0 to -1) := (others => '0');
    variable statevar0 : std_logic_vector(0 to 80) := (others => '0');
    variable state : control_state := STATE0;
    variable nextout : std_logic_vector (0 to 17);
  begin
    if clk'event and clk='1' then
      output <= nextout;
      goto_L5438 := false;
      goto_L5427 := false;
      goto_L5383 := false;
      goto_L5128 := false;
      goto_L5026 := false;
      goto_L4932 := false;
      goto_L4885 := false;
      goto_L4703 := false;
      goto_L4521 := false;
      goto_L4422 := false;
      goto_L4285 := false;
      goto_L4091 := false;
      goto_L4004 := false;
      goto_L3943 := false;
      goto_L3848 := false;
      goto_L3737 := false;
      goto_L3628 := false;
      goto_L3517 := false;
      goto_L3408 := false;
      goto_L3234 := false;
      goto_L3048 := false;
      goto_L2862 := false;
      goto_L2676 := false;
      goto_L2547 := false;
      goto_L2339 := false;
      goto_L2135 := false;
      goto_L1927 := false;
      goto_L1723 := false;
      goto_L1506 := false;
      goto_L1537 := false;
      goto_L1546 := false;
      goto_L1555 := false;
      goto_L1549 := false;
      goto_L1540 := false;
      goto_L1531 := false;
      goto_L1528 := false;
      goto_L1189 := false;
      goto_L1391 := false;
      goto_L1202 := false;
      goto_L1259 := false;
      goto_L1303 := false;
      goto_L1347 := false;
      goto_L1341 := false;
      goto_L1297 := false;
      goto_L1253 := false;
      goto_L1215 := false;
      goto_L1198 := false;
      goto_L814 := false;
      goto_L1115 := false;
      goto_L882 := false;
      goto_L966 := false;
      goto_L1005 := false;
      goto_L1044 := false;
      goto_L1040 := false;
      goto_L1001 := false;
      goto_L962 := false;
      goto_L927 := false;
      goto_L878 := false;
      goto_L732 := false;
      goto_L705 := false;
      goto_L404 := false;
      goto_L314 := false;
      goto_L279 := false;
      goto_L182 := false;
      goto_L225 := false;
      goto_L323 := false;
      goto_L714 := false;
      goto_L1396 := false;
      goto_L1564 := false;
      goto_L1732 := false;
      goto_L1936 := false;
      goto_L2144 := false;
      goto_L2348 := false;
      goto_L2556 := false;
      goto_L2685 := false;
      goto_L2871 := false;
      goto_L3057 := false;
      goto_L3243 := false;
      goto_L3417 := false;
      goto_L3526 := false;
      goto_L3637 := false;
      goto_L3746 := false;
      goto_L3857 := false;
      goto_L3952 := false;
      goto_L4013 := false;
      goto_L4100 := false;
      goto_L4294 := false;
      goto_L4431 := false;
      goto_L4530 := false;
      goto_L4712 := false;
      goto_L4894 := false;
      goto_L5138 := false;
      goto_L5392 := false;
      goto_L5176 := false;
      goto_L5189 := false;
      goto_L5196 := false;
      goto_L5203 := false;
      goto_L5199 := false;
      goto_L5192 := false;
      goto_L5185 := false;
      goto_L5182 := false;
      goto_L5234 := false;
      goto_L5253 := false;
      goto_L5273 := false;
      goto_L5266 := false;
      goto_L5247 := false;
      goto_L5227 := false;
      goto_L5287 := false;
      goto_L5331 := false;
      goto_L5340 := false;
      goto_L5349 := false;
      goto_L5343 := false;
      goto_L5334 := false;
      goto_L5325 := false;
      goto_L5322 := false;
      goto_L4931 := false;
      goto_L5035 := false;
      goto_L5051 := false;
      goto_L5058 := false;
      goto_L5065 := false;
      goto_L5061 := false;
      goto_L5054 := false;
      goto_L5047 := false;
      goto_L5044 := false;
      goto_L5088 := false;
      goto_L5099 := false;
      goto_L5110 := false;
      goto_L5102 := false;
      goto_L5091 := false;
      goto_L5080 := false;
      goto_L5077 := false;
      goto_L4936 := false;
      goto_L4949 := false;
      goto_L4956 := false;
      goto_L4963 := false;
      goto_L4959 := false;
      goto_L4952 := false;
      goto_L4945 := false;
      goto_L4942 := false;
      goto_L4986 := false;
      goto_L4997 := false;
      goto_L5008 := false;
      goto_L5000 := false;
      goto_L4989 := false;
      goto_L4978 := false;
      goto_L4975 := false;
      goto_L4750 := false;
      goto_L4763 := false;
      goto_L4770 := false;
      goto_L4777 := false;
      goto_L4773 := false;
      goto_L4766 := false;
      goto_L4759 := false;
      goto_L4756 := false;
      goto_L4833 := false;
      goto_L4842 := false;
      goto_L4851 := false;
      goto_L4845 := false;
      goto_L4836 := false;
      goto_L4827 := false;
      goto_L4824 := false;
      goto_L4568 := false;
      goto_L4581 := false;
      goto_L4588 := false;
      goto_L4595 := false;
      goto_L4591 := false;
      goto_L4584 := false;
      goto_L4577 := false;
      goto_L4574 := false;
      goto_L4651 := false;
      goto_L4660 := false;
      goto_L4669 := false;
      goto_L4663 := false;
      goto_L4654 := false;
      goto_L4645 := false;
      goto_L4642 := false;
      goto_L4469 := false;
      goto_L4484 := false;
      goto_L4494 := false;
      goto_L4504 := false;
      goto_L4497 := false;
      goto_L4487 := false;
      goto_L4477 := false;
      goto_L4474 := false;
      goto_L4332 := false;
      goto_L4345 := false;
      goto_L4352 := false;
      goto_L4359 := false;
      goto_L4355 := false;
      goto_L4348 := false;
      goto_L4341 := false;
      goto_L4338 := false;
      goto_L4382 := false;
      goto_L4393 := false;
      goto_L4404 := false;
      goto_L4396 := false;
      goto_L4385 := false;
      goto_L4374 := false;
      goto_L4371 := false;
      goto_L4138 := false;
      goto_L4051 := false;
      goto_L3990 := false;
      goto_L3895 := false;
      goto_L3908 := false;
      goto_L3915 := false;
      goto_L3922 := false;
      goto_L3918 := false;
      goto_L3911 := false;
      goto_L3904 := false;
      goto_L3901 := false;
      goto_L3784 := false;
      goto_L3836 := false;
      goto_L3795 := false;
      goto_L3808 := false;
      goto_L3815 := false;
      goto_L3822 := false;
      goto_L3818 := false;
      goto_L3811 := false;
      goto_L3804 := false;
      goto_L3801 := false;
      goto_L3791 := false;
      goto_L3675 := false;
      goto_L3725 := false;
      goto_L3684 := false;
      goto_L3697 := false;
      goto_L3704 := false;
      goto_L3711 := false;
      goto_L3707 := false;
      goto_L3700 := false;
      goto_L3693 := false;
      goto_L3690 := false;
      goto_L3680 := false;
      goto_L3564 := false;
      goto_L3616 := false;
      goto_L3575 := false;
      goto_L3588 := false;
      goto_L3595 := false;
      goto_L3602 := false;
      goto_L3598 := false;
      goto_L3591 := false;
      goto_L3584 := false;
      goto_L3581 := false;
      goto_L3571 := false;
      goto_L3455 := false;
      goto_L3505 := false;
      goto_L3464 := false;
      goto_L3477 := false;
      goto_L3484 := false;
      goto_L3491 := false;
      goto_L3487 := false;
      goto_L3480 := false;
      goto_L3473 := false;
      goto_L3470 := false;
      goto_L3460 := false;
      goto_L3281 := false;
      goto_L3294 := false;
      goto_L3301 := false;
      goto_L3308 := false;
      goto_L3304 := false;
      goto_L3297 := false;
      goto_L3290 := false;
      goto_L3287 := false;
      goto_L3328 := false;
      goto_L3335 := false;
      goto_L3342 := false;
      goto_L3338 := false;
      goto_L3331 := false;
      goto_L3324 := false;
      goto_L3321 := false;
      goto_L3095 := false;
      goto_L3108 := false;
      goto_L3115 := false;
      goto_L3122 := false;
      goto_L3118 := false;
      goto_L3111 := false;
      goto_L3104 := false;
      goto_L3101 := false;
      goto_L3142 := false;
      goto_L3149 := false;
      goto_L3156 := false;
      goto_L3152 := false;
      goto_L3145 := false;
      goto_L3138 := false;
      goto_L3135 := false;
      goto_L3181 := false;
      goto_L3190 := false;
      goto_L3199 := false;
      goto_L3193 := false;
      goto_L3184 := false;
      goto_L3175 := false;
      goto_L3172 := false;
      goto_L2909 := false;
      goto_L2922 := false;
      goto_L2929 := false;
      goto_L2936 := false;
      goto_L2932 := false;
      goto_L2925 := false;
      goto_L2918 := false;
      goto_L2915 := false;
      goto_L2956 := false;
      goto_L2963 := false;
      goto_L2970 := false;
      goto_L2966 := false;
      goto_L2959 := false;
      goto_L2952 := false;
      goto_L2949 := false;
      goto_L2995 := false;
      goto_L3004 := false;
      goto_L3013 := false;
      goto_L3007 := false;
      goto_L2998 := false;
      goto_L2989 := false;
      goto_L2986 := false;
      goto_L2723 := false;
      goto_L2736 := false;
      goto_L2743 := false;
      goto_L2750 := false;
      goto_L2746 := false;
      goto_L2739 := false;
      goto_L2732 := false;
      goto_L2729 := false;
      goto_L2770 := false;
      goto_L2777 := false;
      goto_L2784 := false;
      goto_L2780 := false;
      goto_L2773 := false;
      goto_L2766 := false;
      goto_L2763 := false;
      goto_L2809 := false;
      goto_L2818 := false;
      goto_L2827 := false;
      goto_L2821 := false;
      goto_L2812 := false;
      goto_L2803 := false;
      goto_L2800 := false;
      goto_L2594 := false;
      goto_L2607 := false;
      goto_L2614 := false;
      goto_L2621 := false;
      goto_L2617 := false;
      goto_L2610 := false;
      goto_L2603 := false;
      goto_L2600 := false;
      goto_L2642 := false;
      goto_L2651 := false;
      goto_L2660 := false;
      goto_L2654 := false;
      goto_L2645 := false;
      goto_L2636 := false;
      goto_L2633 := false;
      goto_L2386 := false;
      goto_L2399 := false;
      goto_L2406 := false;
      goto_L2413 := false;
      goto_L2409 := false;
      goto_L2402 := false;
      goto_L2395 := false;
      goto_L2392 := false;
      goto_L2433 := false;
      goto_L2440 := false;
      goto_L2447 := false;
      goto_L2443 := false;
      goto_L2436 := false;
      goto_L2429 := false;
      goto_L2426 := false;
      goto_L2513 := false;
      goto_L2522 := false;
      goto_L2531 := false;
      goto_L2525 := false;
      goto_L2516 := false;
      goto_L2507 := false;
      goto_L2504 := false;
      goto_L2182 := false;
      goto_L2195 := false;
      goto_L2202 := false;
      goto_L2209 := false;
      goto_L2205 := false;
      goto_L2198 := false;
      goto_L2191 := false;
      goto_L2188 := false;
      goto_L2229 := false;
      goto_L2236 := false;
      goto_L2243 := false;
      goto_L2239 := false;
      goto_L2232 := false;
      goto_L2225 := false;
      goto_L2222 := false;
      goto_L2305 := false;
      goto_L2314 := false;
      goto_L2323 := false;
      goto_L2317 := false;
      goto_L2308 := false;
      goto_L2299 := false;
      goto_L2296 := false;
      goto_L1974 := false;
      goto_L1987 := false;
      goto_L1994 := false;
      goto_L2001 := false;
      goto_L1997 := false;
      goto_L1990 := false;
      goto_L1983 := false;
      goto_L1980 := false;
      goto_L2021 := false;
      goto_L2028 := false;
      goto_L2035 := false;
      goto_L2031 := false;
      goto_L2024 := false;
      goto_L2017 := false;
      goto_L2014 := false;
      goto_L2101 := false;
      goto_L2110 := false;
      goto_L2119 := false;
      goto_L2113 := false;
      goto_L2104 := false;
      goto_L2095 := false;
      goto_L2092 := false;
      goto_L1770 := false;
      goto_L1783 := false;
      goto_L1790 := false;
      goto_L1797 := false;
      goto_L1793 := false;
      goto_L1786 := false;
      goto_L1779 := false;
      goto_L1776 := false;
      goto_L1817 := false;
      goto_L1824 := false;
      goto_L1831 := false;
      goto_L1827 := false;
      goto_L1820 := false;
      goto_L1813 := false;
      goto_L1810 := false;
      goto_L1893 := false;
      goto_L1902 := false;
      goto_L1911 := false;
      goto_L1905 := false;
      goto_L1896 := false;
      goto_L1887 := false;
      goto_L1884 := false;
      goto_L1602 := false;
      goto_L1615 := false;
      goto_L1622 := false;
      goto_L1629 := false;
      goto_L1625 := false;
      goto_L1618 := false;
      goto_L1611 := false;
      goto_L1608 := false;
      goto_L1649 := false;
      goto_L1656 := false;
      goto_L1663 := false;
      goto_L1659 := false;
      goto_L1652 := false;
      goto_L1645 := false;
      goto_L1642 := false;
      goto_L1434 := false;
      goto_L1447 := false;
      goto_L1454 := false;
      goto_L1461 := false;
      goto_L1457 := false;
      goto_L1450 := false;
      goto_L1443 := false;
      goto_L1440 := false;
      goto_L770 := false;
      goto_L418 := false;
      goto_L283 := false;
      goto_L0 := false;
      goto_L5439 := false;
      null; -- label L5438
      -- ENTER
      goto_L0 := (state = STATE0);
      if (NOT goto_L0) then
        goto_L182 := (state = STATE182);
        if (NOT goto_L182) then
          goto_L314 := (state = STATE314);
          if (NOT goto_L314) then
            goto_L705 := (state = STATE705);
            if (NOT goto_L705) then
              goto_L814 := (state = STATE814);
              if (NOT goto_L814) then
                goto_L1189 := (state = STATE1189);
                if (NOT goto_L1189) then
                  goto_L1506 := (state = STATE1506);
                  if (NOT goto_L1506) then
                    goto_L1723 := (state = STATE1723);
                    if (NOT goto_L1723) then
                      goto_L1927 := (state = STATE1927);
                      if (NOT goto_L1927) then
                        goto_L2135 := (state = STATE2135);
                        if (NOT goto_L2135) then
                          goto_L2339 := (state = STATE2339);
                          if (NOT goto_L2339) then
                            goto_L2547 := (state = STATE2547);
                            if (NOT goto_L2547) then
                              goto_L2676 := (state = STATE2676);
                              if (NOT goto_L2676) then
                                goto_L2862 := (state = STATE2862);
                                if (NOT goto_L2862) then
                                  goto_L3048 := (state = STATE3048);
                                  if (NOT goto_L3048) then
                                    goto_L3234 := (state = STATE3234);
                                    if (NOT goto_L3234) then
                                      goto_L3408 := (state = STATE3408);
                                      if (NOT goto_L3408) then
                                        goto_L3517 := (state = STATE3517);
                                        if (NOT goto_L3517) then
                                          goto_L3628 := (state = STATE3628);
                                          if (NOT goto_L3628) then
                                            goto_L3737 := (state = STATE3737);
                                            if (NOT goto_L3737) then
                                              goto_L3848 := (state = STATE3848);
                                              if (NOT goto_L3848) then
                                                goto_L3943 := (state = STATE3943);
                                                if (NOT goto_L3943) then
                                                  goto_L4004 := (state = STATE4004);
                                                  if (NOT goto_L4004) then
                                                    goto_L4091 := (state = STATE4091);
                                                    if (NOT goto_L4091) then
                                                      goto_L4285 := (state = STATE4285);
                                                      if (NOT goto_L4285) then
                                                        goto_L4422 := (state = STATE4422);
                                                        if (NOT goto_L4422) then
                                                          goto_L4521 := (state = STATE4521);
                                                          if (NOT goto_L4521) then
                                                            goto_L4703 := (state = STATE4703);
                                                            if (NOT goto_L4703) then
                                                              goto_L4885 := (state = STATE4885);
                                                              if (NOT goto_L4885) then
                                                                goto_L5026 := (state = STATE5026);
                                                                if (NOT goto_L5026) then
                                                                  goto_L5128 := (state = STATE5128);
                                                                  if (NOT goto_L5128) then
                                                                    goto_L5383 := (state = STATE5383);
                                                                    if (NOT goto_L5383) then
                                                                      goto_L5427 := (state = STATE5427);
                                                                      null; -- label L5427
                                                                      r5426 := input;
                                                                      r5428 := statevar0;
                                                                      -- got s@N0 in r5428
                                                                      -- got i@MV in r5426
                                                                      r5432 := rewire_setInputs_185(r5428,r5426);
                                                                      statevar0 := r5432;
                                                                      null;
                                                                      goto_L732 := true;
                                                                    end if;
                                                                    goto_L732 := goto_L732;
                                                                    if (NOT goto_L732) then
                                                                      null; -- label L5383
                                                                      r5382 := input;
                                                                      r5384 := statevar0;
                                                                      -- got s@MM in r5384
                                                                      -- got i@ML in r5382
                                                                      r5388 := rewire_setInputs_185(r5384,r5382);
                                                                      statevar0 := r5388;
                                                                      null;
                                                                      goto_L732 := true;
                                                                    end if;
                                                                    goto_L732 := goto_L732;
                                                                  end if;
                                                                  goto_L732 := goto_L732;
                                                                  if (NOT goto_L732) then
                                                                    null; -- label L5128
                                                                    r5127 := input;
                                                                    r5129 := statevar0;
                                                                    -- got s@M1 in r5129
                                                                    -- got i@M0 in r5127
                                                                    r5133 := rewire_setInputs_185(r5129,r5127);
                                                                    statevar0 := r5133;
                                                                    null;
                                                                    goto_L4932 := true;
                                                                  end if;
                                                                  goto_L4932 := goto_L4932;
                                                                end if;
                                                                goto_L4932 := goto_L4932;
                                                                if (NOT goto_L4932) then
                                                                  goto_L732 := goto_L732;
                                                                  if (NOT goto_L732) then
                                                                    null; -- label L5026
                                                                    r5025 := input;
                                                                    r5027 := statevar0;
                                                                    -- got s@LP in r5027
                                                                    -- got i@LO in r5025
                                                                    r5031 := rewire_setInputs_185(r5027,r5025);
                                                                    statevar0 := r5031;
                                                                    null;
                                                                    goto_L4932 := true;
                                                                  end if;
                                                                  goto_L4932 := goto_L4932;
                                                                end if;
                                                                goto_L4932 := goto_L4932;
                                                                if (NOT goto_L4932) then
                                                                  goto_L732 := goto_L732;
                                                                end if;
                                                                goto_L732 := goto_L732;
                                                                if (NOT goto_L732) then
                                                                  null; -- label L4932
                                                                  -- end case
                                                                  null;
                                                                  goto_L732 := true;
                                                                end if;
                                                                goto_L732 := goto_L732;
                                                              end if;
                                                              goto_L732 := goto_L732;
                                                              if (NOT goto_L732) then
                                                                null; -- label L4885
                                                                r4884 := input;
                                                                r4886 := statevar0;
                                                                -- got s@LE in r4886
                                                                -- got i@LD in r4884
                                                                r4890 := rewire_setInputs_185(r4886,r4884);
                                                                statevar0 := r4890;
                                                                null;
                                                                goto_L732 := true;
                                                              end if;
                                                              goto_L732 := goto_L732;
                                                            end if;
                                                            goto_L732 := goto_L732;
                                                            if (NOT goto_L732) then
                                                              null; -- label L4703
                                                              r4702 := input;
                                                              r4704 := statevar0;
                                                              -- got s@KR in r4704
                                                              -- got i@KQ in r4702
                                                              r4708 := rewire_setInputs_185(r4704,r4702);
                                                              statevar0 := r4708;
                                                              null;
                                                              goto_L732 := true;
                                                            end if;
                                                            goto_L732 := goto_L732;
                                                          end if;
                                                          goto_L732 := goto_L732;
                                                          if (NOT goto_L732) then
                                                            null; -- label L4521
                                                            r4520 := input;
                                                            r4522 := statevar0;
                                                            -- got s@K8 in r4522
                                                            -- got i@K7 in r4520
                                                            r4526 := rewire_setInputs_185(r4522,r4520);
                                                            statevar0 := r4526;
                                                            null;
                                                            goto_L732 := true;
                                                          end if;
                                                          goto_L732 := goto_L732;
                                                        end if;
                                                        goto_L732 := goto_L732;
                                                        if (NOT goto_L732) then
                                                          null; -- label L4422
                                                          r4421 := input;
                                                          r4423 := statevar0;
                                                          -- got s@K0 in r4423
                                                          -- got i@JV in r4421
                                                          r4427 := rewire_setInputs_185(r4423,r4421);
                                                          statevar0 := r4427;
                                                          null;
                                                          goto_L732 := true;
                                                        end if;
                                                        goto_L732 := goto_L732;
                                                      end if;
                                                      goto_L732 := goto_L732;
                                                      if (NOT goto_L732) then
                                                        null; -- label L4285
                                                        r4284 := input;
                                                        r4286 := statevar0;
                                                        -- got s@JM in r4286
                                                        -- got i@JL in r4284
                                                        r4290 := rewire_setInputs_185(r4286,r4284);
                                                        statevar0 := r4290;
                                                        null;
                                                        goto_L732 := true;
                                                      end if;
                                                      goto_L732 := goto_L732;
                                                    end if;
                                                    goto_L732 := goto_L732;
                                                    if (NOT goto_L732) then
                                                      null; -- label L4091
                                                      r4090 := input;
                                                      r4092 := statevar0;
                                                      -- got s@J4 in r4092
                                                      -- got i@J3 in r4090
                                                      r4096 := rewire_setInputs_185(r4092,r4090);
                                                      statevar0 := r4096;
                                                      null;
                                                      goto_L732 := true;
                                                    end if;
                                                    goto_L732 := goto_L732;
                                                  end if;
                                                  goto_L732 := goto_L732;
                                                  if (NOT goto_L732) then
                                                    null; -- label L4004
                                                    r4003 := input;
                                                    r4005 := statevar0;
                                                    -- got s@IS in r4005
                                                    -- got i@IR in r4003
                                                    r4009 := rewire_setInputs_185(r4005,r4003);
                                                    statevar0 := r4009;
                                                    null;
                                                    goto_L732 := true;
                                                  end if;
                                                  goto_L732 := goto_L732;
                                                end if;
                                                goto_L732 := goto_L732;
                                                if (NOT goto_L732) then
                                                  null; -- label L3943
                                                  r3942 := input;
                                                  r3944 := statevar0;
                                                  -- got s@IL in r3944
                                                  -- got i@IK in r3942
                                                  r3948 := rewire_setInputs_185(r3944,r3942);
                                                  statevar0 := r3948;
                                                  null;
                                                  goto_L732 := true;
                                                end if;
                                                goto_L732 := goto_L732;
                                              end if;
                                              goto_L732 := goto_L732;
                                              if (NOT goto_L732) then
                                                null; -- label L3848
                                                r3847 := input;
                                                r3849 := statevar0;
                                                -- got s@IB in r3849
                                                -- got i@IA in r3847
                                                r3853 := rewire_setInputs_185(r3849,r3847);
                                                statevar0 := r3853;
                                                null;
                                                goto_L732 := true;
                                              end if;
                                              goto_L732 := goto_L732;
                                            end if;
                                            goto_L732 := goto_L732;
                                            if (NOT goto_L732) then
                                              null; -- label L3737
                                              r3736 := input;
                                              r3738 := statevar0;
                                              -- got s@HV in r3738
                                              -- got i@HU in r3736
                                              r3742 := rewire_setInputs_185(r3738,r3736);
                                              statevar0 := r3742;
                                              null;
                                              goto_L732 := true;
                                            end if;
                                            goto_L732 := goto_L732;
                                          end if;
                                          goto_L732 := goto_L732;
                                          if (NOT goto_L732) then
                                            null; -- label L3628
                                            r3627 := input;
                                            r3629 := statevar0;
                                            -- got s@HJ in r3629
                                            -- got i@HI in r3627
                                            r3633 := rewire_setInputs_185(r3629,r3627);
                                            statevar0 := r3633;
                                            null;
                                            goto_L732 := true;
                                          end if;
                                          goto_L732 := goto_L732;
                                        end if;
                                        goto_L732 := goto_L732;
                                        if (NOT goto_L732) then
                                          null; -- label L3517
                                          r3516 := input;
                                          r3518 := statevar0;
                                          -- got s@H7 in r3518
                                          -- got i@H6 in r3516
                                          r3522 := rewire_setInputs_185(r3518,r3516);
                                          statevar0 := r3522;
                                          null;
                                          goto_L732 := true;
                                        end if;
                                        goto_L732 := goto_L732;
                                      end if;
                                      goto_L732 := goto_L732;
                                      if (NOT goto_L732) then
                                        null; -- label L3408
                                        r3407 := input;
                                        r3409 := statevar0;
                                        -- got s@GR in r3409
                                        -- got i@GQ in r3407
                                        r3413 := rewire_setInputs_185(r3409,r3407);
                                        statevar0 := r3413;
                                        null;
                                        goto_L732 := true;
                                      end if;
                                      goto_L732 := goto_L732;
                                    end if;
                                    goto_L732 := goto_L732;
                                    if (NOT goto_L732) then
                                      null; -- label L3234
                                      r3233 := input;
                                      r3235 := statevar0;
                                      -- got s@G6 in r3235
                                      -- got i@G5 in r3233
                                      r3239 := rewire_setInputs_185(r3235,r3233);
                                      statevar0 := r3239;
                                      null;
                                      goto_L732 := true;
                                    end if;
                                    goto_L732 := goto_L732;
                                  end if;
                                  goto_L732 := goto_L732;
                                  if (NOT goto_L732) then
                                    null; -- label L3048
                                    r3047 := input;
                                    r3049 := statevar0;
                                    -- got s@FJ in r3049
                                    -- got i@FI in r3047
                                    r3053 := rewire_setInputs_185(r3049,r3047);
                                    statevar0 := r3053;
                                    null;
                                    goto_L732 := true;
                                  end if;
                                  goto_L732 := goto_L732;
                                end if;
                                goto_L732 := goto_L732;
                                if (NOT goto_L732) then
                                  null; -- label L2862
                                  r2861 := input;
                                  r2863 := statevar0;
                                  -- got s@F0 in r2863
                                  -- got i@EV in r2861
                                  r2867 := rewire_setInputs_185(r2863,r2861);
                                  statevar0 := r2867;
                                  null;
                                  goto_L732 := true;
                                end if;
                                goto_L732 := goto_L732;
                              end if;
                              goto_L732 := goto_L732;
                              if (NOT goto_L732) then
                                null; -- label L2676
                                r2675 := input;
                                r2677 := statevar0;
                                -- got s@ED in r2677
                                -- got i@EC in r2675
                                r2681 := rewire_setInputs_185(r2677,r2675);
                                statevar0 := r2681;
                                null;
                                goto_L732 := true;
                              end if;
                              goto_L732 := goto_L732;
                            end if;
                            goto_L732 := goto_L732;
                            if (NOT goto_L732) then
                              null; -- label L2547
                              r2546 := input;
                              r2548 := statevar0;
                              -- got s@E1 in r2548
                              -- got i@E0 in r2546
                              r2552 := rewire_setInputs_185(r2548,r2546);
                              statevar0 := r2552;
                              null;
                              goto_L732 := true;
                            end if;
                            goto_L732 := goto_L732;
                          end if;
                          goto_L732 := goto_L732;
                          if (NOT goto_L732) then
                            null; -- label L2339
                            r2338 := input;
                            r2340 := statevar0;
                            -- got s@DA in r2340
                            -- got i@D9 in r2338
                            r2344 := rewire_setInputs_185(r2340,r2338);
                            statevar0 := r2344;
                            null;
                            goto_L732 := true;
                          end if;
                          goto_L732 := goto_L732;
                        end if;
                        goto_L732 := goto_L732;
                        if (NOT goto_L732) then
                          null; -- label L2135
                          r2134 := input;
                          r2136 := statevar0;
                          -- got s@CL in r2136
                          -- got i@CK in r2134
                          r2140 := rewire_setInputs_185(r2136,r2134);
                          statevar0 := r2140;
                          null;
                          goto_L732 := true;
                        end if;
                        goto_L732 := goto_L732;
                      end if;
                      goto_L732 := goto_L732;
                      if (NOT goto_L732) then
                        null; -- label L1927
                        r1926 := input;
                        r1928 := statevar0;
                        -- got s@BU in r1928
                        -- got i@BT in r1926
                        r1932 := rewire_setInputs_185(r1928,r1926);
                        statevar0 := r1932;
                        null;
                        goto_L732 := true;
                      end if;
                      goto_L732 := goto_L732;
                    end if;
                    goto_L732 := goto_L732;
                    if (NOT goto_L732) then
                      null; -- label L1723
                      r1722 := input;
                      r1724 := statevar0;
                      -- got s@B9 in r1724
                      -- got i@B8 in r1722
                      r1728 := rewire_setInputs_185(r1724,r1722);
                      statevar0 := r1728;
                      null;
                      goto_L732 := true;
                    end if;
                    goto_L732 := goto_L732;
                  end if;
                  goto_L732 := goto_L732;
                  if (NOT goto_L732) then
                    null; -- label L1506
                    r1505 := input;
                    r1507 := statevar0;
                    -- got s@AC in r1507
                    -- got i@AB in r1505
                    r1511 := rewire_setInputs_185(r1507,r1505);
                    statevar0 := r1511;
                    r1514 := statevar0;
                    -- got s@AE in r1514
                    r1517 := rewire_inputs_229(r1514);
                    -- got i@AF in r1517
                    r1520 := rewire_dataIn_717(r1517);
                    r1522 := statevar0;
                    -- got b0@9R in r1407
                    -- got b1@9S in r1409
                    r1526 := rewire_mkReg_883(r1407,r1409);
                    b1529 := ("00" = r1526(0 to 1));
                    goto_L1531 := b1529;
                    if (NOT goto_L1531) then
                      goto_L1537 := (NOT b1529);
                      null; -- label L1537
                      -- alt exit (no match)
                      b1538 := ("01" = r1526(0 to 1));
                      goto_L1540 := b1538;
                      if (NOT goto_L1540) then
                        goto_L1546 := (NOT b1538);
                        null; -- label L1546
                        -- alt exit (no match)
                        b1547 := ("10" = r1526(0 to 1));
                        goto_L1549 := b1547;
                        if (NOT goto_L1549) then
                          goto_L1555 := (NOT b1547);
                          null; -- label L1555
                          -- alt exit (no match)
                          -- final pat
                          -- got s@AH in r1522
                          -- got v@AG in r1520
                          r1559 := rewire_setR3_1349(r1522,r1520);
                          statevar0 := r1559;
                          null;
                          goto_L1528 := true;
                        end if;
                        goto_L1528 := goto_L1528;
                        if (NOT goto_L1528) then
                          null; -- label L1549
                          -- got s@AH in r1522
                          -- got v@AG in r1520
                          r1551 := rewire_setR2_1306(r1522,r1520);
                          statevar0 := r1551;
                          null;
                          goto_L1528 := true;
                        end if;
                        goto_L1528 := goto_L1528;
                      end if;
                      goto_L1528 := goto_L1528;
                      if (NOT goto_L1528) then
                        null; -- label L1540
                        -- got s@AH in r1522
                        -- got v@AG in r1520
                        r1542 := rewire_setR1_1262(r1522,r1520);
                        statevar0 := r1542;
                        null;
                        goto_L1528 := true;
                      end if;
                      goto_L1528 := goto_L1528;
                    end if;
                    goto_L1528 := goto_L1528;
                    if (NOT goto_L1528) then
                      null; -- label L1531
                      -- got s@AH in r1522
                      -- got v@AG in r1520
                      r1533 := rewire_setR0_1218(r1522,r1520);
                      statevar0 := r1533;
                      null;
                      goto_L1528 := true;
                    end if;
                    goto_L1528 := goto_L1528;
                    null; -- label L1528
                    -- end case
                    null;
                    goto_L732 := true;
                  end if;
                  goto_L732 := goto_L732;
                end if;
                goto_L732 := goto_L732;
                if (NOT goto_L732) then
                  null; -- label L1189
                  r1188 := input;
                  r1190 := statevar0;
                  -- got s@9L in r1190
                  -- got i@9K in r1188
                  r1194 := rewire_setInputs_185(r1190,r1188);
                  statevar0 := r1194;
                  -- got rEn@8D in r743
                  b1199 := ("1" = r743(0 to 0));
                  goto_L1202 := b1199;
                  if (NOT goto_L1202) then
                    goto_L1391 := (NOT b1199);
                    null; -- label L1391
                    -- alt exit (no match)
                    -- final pat
                    null;
                    null;
                    goto_L1198 := true;
                  end if;
                  goto_L1198 := goto_L1198;
                  if (NOT goto_L1198) then
                    null; -- label L1202
                    r1201 := statevar0;
                    -- got s@9N in r1201
                    r1204 := rewire_inputs_229(r1201);
                    -- got i@9O in r1204
                    r1207 := rewire_dataIn_717(r1204);
                    r1209 := statevar0;
                    -- got b0@8F in r747
                    -- got b1@8G in r749
                    r1213 := rewire_mkReg_883(r747,r749);
                    b1216 := ("00" = r1213(0 to 1));
                    goto_L1253 := b1216;
                    if (NOT goto_L1253) then
                      goto_L1259 := (NOT b1216);
                      null; -- label L1259
                      -- alt exit (no match)
                      b1260 := ("01" = r1213(0 to 1));
                      goto_L1297 := b1260;
                      if (NOT goto_L1297) then
                        goto_L1303 := (NOT b1260);
                        null; -- label L1303
                        -- alt exit (no match)
                        b1304 := ("10" = r1213(0 to 1));
                        goto_L1341 := b1304;
                        if (NOT goto_L1341) then
                          goto_L1347 := (NOT b1304);
                          null; -- label L1347
                          -- alt exit (no match)
                          -- final pat
                          -- got s@9Q in r1209
                          -- got v@9P in r1207
                          r1386 := rewire_setR3_1349(r1209,r1207);
                          statevar0 := r1386;
                          null;
                          goto_L1215 := true;
                        end if;
                        goto_L1215 := goto_L1215;
                        if (NOT goto_L1215) then
                          null; -- label L1341
                          -- got s@9Q in r1209
                          -- got v@9P in r1207
                          r1343 := rewire_setR2_1306(r1209,r1207);
                          statevar0 := r1343;
                          null;
                          goto_L1215 := true;
                        end if;
                        goto_L1215 := goto_L1215;
                      end if;
                      goto_L1215 := goto_L1215;
                      if (NOT goto_L1215) then
                        null; -- label L1297
                        -- got s@9Q in r1209
                        -- got v@9P in r1207
                        r1299 := rewire_setR1_1262(r1209,r1207);
                        statevar0 := r1299;
                        null;
                        goto_L1215 := true;
                      end if;
                      goto_L1215 := goto_L1215;
                    end if;
                    goto_L1215 := goto_L1215;
                    if (NOT goto_L1215) then
                      null; -- label L1253
                      -- got s@9Q in r1209
                      -- got v@9P in r1207
                      r1255 := rewire_setR0_1218(r1209,r1207);
                      statevar0 := r1255;
                      null;
                      goto_L1215 := true;
                    end if;
                    goto_L1215 := goto_L1215;
                    null; -- label L1215
                    -- end case
                    null;
                    goto_L1198 := true;
                  end if;
                  goto_L1198 := goto_L1198;
                  null; -- label L1198
                  -- end case
                  null;
                  goto_L732 := true;
                end if;
                goto_L732 := goto_L732;
              end if;
              goto_L732 := goto_L732;
              if (NOT goto_L732) then
                null; -- label L814
                r813 := input;
                r815 := statevar0;
                -- got s@8Q in r815
                -- got i@8P in r813
                r819 := rewire_setInputs_185(r815,r813);
                statevar0 := r819;
                r822 := statevar0;
                -- got s@8S in r822
                r825 := rewire_inputs_229(r822);
                -- got i@8T in r825
                r828 := rewire_dataIn_717(r825);
                r830 := statevar0;
                -- got s@8V in r830
                r833 := rewire_outputs_144(r830);
                r835 := statevar0;
                -- got s@91 in r835
                -- got o@90 in r833
                -- got a@8U in r828
                r840 := rewire_setAddrOut_782(r833,r828);
                r842 := rewire_setOutputs_91(r835,r840);
                statevar0 := r842;
                r845 := statevar0;
                -- got s@93 in r845
                r848 := rewire_outputs_144(r845);
                r850 := statevar0;
                -- got s@95 in r850
                -- got o@94 in r848
                -- got wEn@8E in r745
                r872 := rewire_setWeOut_853(r848,r745);
                r874 := rewire_setOutputs_91(r850,r872);
                statevar0 := r874;
                -- got wEn@8E in r745
                b879 := ("1" = r745(0 to 0));
                goto_L882 := b879;
                if (NOT goto_L882) then
                  goto_L1115 := (NOT b879);
                  null; -- label L1115
                  -- alt exit (no match)
                  -- final pat
                  null;
                  null;
                  goto_L878 := true;
                end if;
                goto_L878 := goto_L878;
                if (NOT goto_L878) then
                  null; -- label L882
                  r881 := statevar0;
                  -- got b0@8F in r747
                  -- got b1@8G in r749
                  r924 := rewire_mkReg_883(r747,r749);
                  b928 := ("00" = r924(0 to 1));
                  goto_L962 := b928;
                  if (NOT goto_L962) then
                    goto_L966 := (NOT b928);
                    null; -- label L966
                    -- alt exit (no match)
                    b967 := ("01" = r924(0 to 1));
                    goto_L1001 := b967;
                    if (NOT goto_L1001) then
                      goto_L1005 := (NOT b967);
                      null; -- label L1005
                      -- alt exit (no match)
                      b1006 := ("10" = r924(0 to 1));
                      goto_L1040 := b1006;
                      if (NOT goto_L1040) then
                        goto_L1044 := (NOT b1006);
                        null; -- label L1044
                        -- alt exit (no match)
                        -- final pat
                        -- got s@97 in r881
                        r1079 := rewire_r3_1046(r881);
                        r926 := r1079;
                        goto_L927 := true;
                      end if;
                      goto_L927 := goto_L927;
                      if (NOT goto_L927) then
                        null; -- label L1040
                        -- got s@97 in r881
                        r1041 := rewire_r2_1008(r881);
                        r926 := r1041;
                        goto_L927 := true;
                      end if;
                      goto_L927 := goto_L927;
                    end if;
                    goto_L927 := goto_L927;
                    if (NOT goto_L927) then
                      null; -- label L1001
                      -- got s@97 in r881
                      r1002 := rewire_r1_969(r881);
                      r926 := r1002;
                      goto_L927 := true;
                    end if;
                    goto_L927 := goto_L927;
                  end if;
                  goto_L927 := goto_L927;
                  if (NOT goto_L927) then
                    null; -- label L962
                    -- got s@97 in r881
                    r963 := rewire_r0_930(r881);
                    r926 := r963;
                    goto_L927 := true;
                  end if;
                  goto_L927 := goto_L927;
                  null; -- label L927
                  -- end case
                  r1082 := statevar0;
                  -- got s@99 in r1082
                  r1085 := rewire_outputs_144(r1082);
                  r1087 := statevar0;
                  -- got s@9B in r1087
                  -- got o@9A in r1085
                  -- got d@98 in r926
                  r1109 := rewire_setDataOut_1090(r1085,r926);
                  r1111 := rewire_setOutputs_91(r1087,r1109);
                  statevar0 := r1111;
                  null;
                  goto_L878 := true;
                end if;
                goto_L878 := goto_L878;
                null; -- label L878
                -- end case
                r1119 := statevar0;
                -- got pc@8I in r772
                r1122 := statevar0;
                -- got s@9F in r1122
                -- got pc'@9E in r772
                r1161 := oneW8;
                r1163 := plusW8(r772,r1161);
                -- final pat
                r1167 := r1163(0 to 0);
                r1169 := r1163(1 to 8);
                b1171 := true;
                b1173 := true;
                -- got x@9G in r1169
                r1165 := r1169;
                -- end case
                r1178 := rewire_setPC_1124(r1122,r1165);
                statevar0 := r1178;
                r1181 := statevar0;
                -- got s@9I in r1181
                r1184 := rewire_outputs_144(r1181);
                -- got o@9J in r1184
                nextout := r1184;
                state := STATE1189;
                goto_L5439 := true;
              end if;
              goto_L5439 := goto_L5439;
              if (NOT goto_L5439) then
                null; -- label L732
                -- end case
                null;
                goto_L404 := true;
              end if;
              goto_L404 := goto_L404;
            end if;
            goto_L404 := goto_L404;
            if (NOT goto_L404) then
              goto_L5439 := goto_L5439;
              if (NOT goto_L5439) then
                null; -- label L705
                r704 := input;
                r706 := statevar0;
                -- got s@8C in r706
                -- got i@8B in r704
                r710 := rewire_setInputs_185(r706,r704);
                statevar0 := r710;
                null;
                goto_L404 := true;
              end if;
              goto_L404 := goto_L404;
            end if;
            goto_L404 := goto_L404;
            if (NOT goto_L404) then
              goto_L5439 := goto_L5439;
            end if;
            goto_L5439 := goto_L5439;
            if (NOT goto_L5439) then
              null; -- label L404
              -- end case
              null;
              goto_L279 := true;
            end if;
            goto_L279 := goto_L279;
          end if;
          goto_L279 := goto_L279;
          if (NOT goto_L279) then
            goto_L5439 := goto_L5439;
            if (NOT goto_L5439) then
              null; -- label L314
              r313 := input;
              r315 := statevar0;
              -- got s@7N in r315
              -- got i@7M in r313
              r319 := rewire_setInputs_185(r315,r313);
              statevar0 := r319;
              null;
              goto_L279 := true;
            end if;
            goto_L279 := goto_L279;
          end if;
          goto_L279 := goto_L279;
          if (NOT goto_L279) then
            goto_L5439 := goto_L5439;
          end if;
          goto_L5439 := goto_L5439;
          if (NOT goto_L5439) then
            null; -- label L279
            -- end case
            goto_L225 := true;
          end if;
          goto_L225 := goto_L225;
        end if;
        goto_L225 := goto_L225;
        if (NOT goto_L225) then
          goto_L5439 := goto_L5439;
          if (NOT goto_L5439) then
            null; -- label L182
            r181 := input;
            r183 := statevar0;
            -- got s@NB in r183
            -- got i@NA in r181
            r222 := rewire_setInputs_185(r183,r181);
            statevar0 := r222;
            goto_L225 := true;
          end if;
          goto_L225 := goto_L225;
        end if;
        goto_L225 := goto_L225;
        if (NOT goto_L225) then
          goto_L5439 := goto_L5439;
        end if;
        goto_L5439 := goto_L5439;
        if (NOT goto_L5439) then
          null; -- label L225
          -- loop in
          r227 := statevar0;
          -- got s@7C in r227
          r262 := rewire_inputs_229(r227);
          -- got inp@7D in r262
          r277 := rewire_rstIn_264(r262);
          b280 := ("1" = r277(0 to 0));
          goto_L283 := b280;
          if (NOT goto_L283) then
            goto_L323 := (NOT b280);
            null; -- label L323
            -- alt exit (no match)
            -- final pat
            r325 := statevar0;
            -- got s@7O in r325
            -- final pat
            r330 := r325(0 to 9);
            r332 := r325(10 to 27);
            r334 := r325(28 to 28);
            r336 := r325(29 to 29);
            r338 := r325(30 to 30);
            r340 := r325(31 to 38);
            r342 := r325(39 to 39);
            r344 := r325(40 to 40);
            r346 := r325(41 to 48);
            r348 := r325(49 to 56);
            r350 := r325(57 to 64);
            r352 := r325(65 to 72);
            r354 := r325(73 to 80);
            b356 := true;
            b358 := true;
            b360 := true;
            b362 := true;
            b364 := true;
            b366 := true;
            b368 := true;
            b370 := true;
            b372 := true;
            b374 := true;
            b376 := true;
            b378 := true;
            b380 := true;
            -- got ie@7P in r338
            r328 := r338;
            -- end case
            null;
            -- got ie@7Q in r328
            -- got inp@7D in r262
            r400 := rewire_intIn_387(r262);
            r402 := (r328 & r400);
            b405 := true;
            r407 := r402(0 to 0);
            r409 := r402(1 to 1);
            b411 := ("1" = r407(0 to 0));
            b413 := ("1" = r409(0 to 0));
            b415 := (b405 AND (b411 AND b413));
            goto_L418 := b415;
            if (NOT goto_L418) then
              goto_L714 := (NOT b415);
              null; -- label L714
              -- alt exit (no match)
              b715 := true;
              -- got inp@7D in r262
              r730 := rewire_dataIn_717(r262);
              b733 := true;
              r735 := r730(0 to 0);
              r737 := r730(1 to 1);
              r739 := r730(2 to 2);
              r741 := r730(3 to 3);
              r743 := r730(4 to 4);
              r745 := r730(5 to 5);
              r747 := r730(6 to 6);
              r749 := r730(7 to 7);
              b751 := ("0" = r735(0 to 0));
              b753 := ("0" = r737(0 to 0));
              b755 := ("0" = r739(0 to 0));
              b757 := ("0" = r741(0 to 0));
              b759 := true;
              b761 := true;
              b763 := true;
              b765 := true;
              b767 := (b733 AND (b751 AND (b753 AND (b755 AND (b757 AND (b759 AND (b761 AND (b763 AND b765))))))));
              goto_L770 := b767;
              if (NOT goto_L770) then
                goto_L1396 := (NOT b767);
                null; -- label L1396
                -- alt exit (no match)
                b1397 := true;
                r1399 := r730(0 to 0);
                r1401 := r730(1 to 1);
                r1403 := r730(2 to 2);
                r1405 := r730(3 to 3);
                r1407 := r730(4 to 4);
                r1409 := r730(5 to 5);
                r1411 := r730(6 to 6);
                r1413 := r730(7 to 7);
                b1415 := ("0" = r1399(0 to 0));
                b1417 := ("0" = r1401(0 to 0));
                b1419 := ("0" = r1403(0 to 0));
                b1421 := ("1" = r1405(0 to 0));
                b1423 := true;
                b1425 := true;
                b1427 := true;
                b1429 := true;
                b1431 := (b1397 AND (b1415 AND (b1417 AND (b1419 AND (b1421 AND (b1423 AND (b1425 AND (b1427 AND b1429))))))));
                goto_L1434 := b1431;
                if (NOT goto_L1434) then
                  goto_L1564 := (NOT b1431);
                  null; -- label L1564
                  -- alt exit (no match)
                  b1565 := true;
                  r1567 := r730(0 to 0);
                  r1569 := r730(1 to 1);
                  r1571 := r730(2 to 2);
                  r1573 := r730(3 to 3);
                  r1575 := r730(4 to 4);
                  r1577 := r730(5 to 5);
                  r1579 := r730(6 to 6);
                  r1581 := r730(7 to 7);
                  b1583 := ("0" = r1567(0 to 0));
                  b1585 := ("0" = r1569(0 to 0));
                  b1587 := ("1" = r1571(0 to 0));
                  b1589 := ("0" = r1573(0 to 0));
                  b1591 := true;
                  b1593 := true;
                  b1595 := true;
                  b1597 := true;
                  b1599 := (b1565 AND (b1583 AND (b1585 AND (b1587 AND (b1589 AND (b1591 AND (b1593 AND (b1595 AND b1597))))))));
                  goto_L1602 := b1599;
                  if (NOT goto_L1602) then
                    goto_L1732 := (NOT b1599);
                    null; -- label L1732
                    -- alt exit (no match)
                    b1733 := true;
                    r1735 := r730(0 to 0);
                    r1737 := r730(1 to 1);
                    r1739 := r730(2 to 2);
                    r1741 := r730(3 to 3);
                    r1743 := r730(4 to 4);
                    r1745 := r730(5 to 5);
                    r1747 := r730(6 to 6);
                    r1749 := r730(7 to 7);
                    b1751 := ("0" = r1735(0 to 0));
                    b1753 := ("0" = r1737(0 to 0));
                    b1755 := ("1" = r1739(0 to 0));
                    b1757 := ("1" = r1741(0 to 0));
                    b1759 := true;
                    b1761 := true;
                    b1763 := true;
                    b1765 := true;
                    b1767 := (b1733 AND (b1751 AND (b1753 AND (b1755 AND (b1757 AND (b1759 AND (b1761 AND (b1763 AND b1765))))))));
                    goto_L1770 := b1767;
                    if (NOT goto_L1770) then
                      goto_L1936 := (NOT b1767);
                      null; -- label L1936
                      -- alt exit (no match)
                      b1937 := true;
                      r1939 := r730(0 to 0);
                      r1941 := r730(1 to 1);
                      r1943 := r730(2 to 2);
                      r1945 := r730(3 to 3);
                      r1947 := r730(4 to 4);
                      r1949 := r730(5 to 5);
                      r1951 := r730(6 to 6);
                      r1953 := r730(7 to 7);
                      b1955 := ("0" = r1939(0 to 0));
                      b1957 := ("1" = r1941(0 to 0));
                      b1959 := ("0" = r1943(0 to 0));
                      b1961 := ("0" = r1945(0 to 0));
                      b1963 := true;
                      b1965 := true;
                      b1967 := true;
                      b1969 := true;
                      b1971 := (b1937 AND (b1955 AND (b1957 AND (b1959 AND (b1961 AND (b1963 AND (b1965 AND (b1967 AND b1969))))))));
                      goto_L1974 := b1971;
                      if (NOT goto_L1974) then
                        goto_L2144 := (NOT b1971);
                        null; -- label L2144
                        -- alt exit (no match)
                        b2145 := true;
                        r2147 := r730(0 to 0);
                        r2149 := r730(1 to 1);
                        r2151 := r730(2 to 2);
                        r2153 := r730(3 to 3);
                        r2155 := r730(4 to 4);
                        r2157 := r730(5 to 5);
                        r2159 := r730(6 to 6);
                        r2161 := r730(7 to 7);
                        b2163 := ("0" = r2147(0 to 0));
                        b2165 := ("1" = r2149(0 to 0));
                        b2167 := ("0" = r2151(0 to 0));
                        b2169 := ("1" = r2153(0 to 0));
                        b2171 := true;
                        b2173 := true;
                        b2175 := true;
                        b2177 := true;
                        b2179 := (b2145 AND (b2163 AND (b2165 AND (b2167 AND (b2169 AND (b2171 AND (b2173 AND (b2175 AND b2177))))))));
                        goto_L2182 := b2179;
                        if (NOT goto_L2182) then
                          goto_L2348 := (NOT b2179);
                          null; -- label L2348
                          -- alt exit (no match)
                          b2349 := true;
                          r2351 := r730(0 to 0);
                          r2353 := r730(1 to 1);
                          r2355 := r730(2 to 2);
                          r2357 := r730(3 to 3);
                          r2359 := r730(4 to 4);
                          r2361 := r730(5 to 5);
                          r2363 := r730(6 to 6);
                          r2365 := r730(7 to 7);
                          b2367 := ("0" = r2351(0 to 0));
                          b2369 := ("1" = r2353(0 to 0));
                          b2371 := ("1" = r2355(0 to 0));
                          b2373 := ("0" = r2357(0 to 0));
                          b2375 := true;
                          b2377 := true;
                          b2379 := true;
                          b2381 := true;
                          b2383 := (b2349 AND (b2367 AND (b2369 AND (b2371 AND (b2373 AND (b2375 AND (b2377 AND (b2379 AND b2381))))))));
                          goto_L2386 := b2383;
                          if (NOT goto_L2386) then
                            goto_L2556 := (NOT b2383);
                            null; -- label L2556
                            -- alt exit (no match)
                            b2557 := true;
                            r2559 := r730(0 to 0);
                            r2561 := r730(1 to 1);
                            r2563 := r730(2 to 2);
                            r2565 := r730(3 to 3);
                            r2567 := r730(4 to 4);
                            r2569 := r730(5 to 5);
                            r2571 := r730(6 to 6);
                            r2573 := r730(7 to 7);
                            b2575 := ("0" = r2559(0 to 0));
                            b2577 := ("1" = r2561(0 to 0));
                            b2579 := ("1" = r2563(0 to 0));
                            b2581 := ("1" = r2565(0 to 0));
                            b2583 := true;
                            b2585 := true;
                            b2587 := true;
                            b2589 := true;
                            b2591 := (b2557 AND (b2575 AND (b2577 AND (b2579 AND (b2581 AND (b2583 AND (b2585 AND (b2587 AND b2589))))))));
                            goto_L2594 := b2591;
                            if (NOT goto_L2594) then
                              goto_L2685 := (NOT b2591);
                              null; -- label L2685
                              -- alt exit (no match)
                              b2686 := true;
                              r2688 := r730(0 to 0);
                              r2690 := r730(1 to 1);
                              r2692 := r730(2 to 2);
                              r2694 := r730(3 to 3);
                              r2696 := r730(4 to 4);
                              r2698 := r730(5 to 5);
                              r2700 := r730(6 to 6);
                              r2702 := r730(7 to 7);
                              b2704 := ("1" = r2688(0 to 0));
                              b2706 := ("0" = r2690(0 to 0));
                              b2708 := ("0" = r2692(0 to 0));
                              b2710 := ("0" = r2694(0 to 0));
                              b2712 := true;
                              b2714 := true;
                              b2716 := true;
                              b2718 := true;
                              b2720 := (b2686 AND (b2704 AND (b2706 AND (b2708 AND (b2710 AND (b2712 AND (b2714 AND (b2716 AND b2718))))))));
                              goto_L2723 := b2720;
                              if (NOT goto_L2723) then
                                goto_L2871 := (NOT b2720);
                                null; -- label L2871
                                -- alt exit (no match)
                                b2872 := true;
                                r2874 := r730(0 to 0);
                                r2876 := r730(1 to 1);
                                r2878 := r730(2 to 2);
                                r2880 := r730(3 to 3);
                                r2882 := r730(4 to 4);
                                r2884 := r730(5 to 5);
                                r2886 := r730(6 to 6);
                                r2888 := r730(7 to 7);
                                b2890 := ("1" = r2874(0 to 0));
                                b2892 := ("0" = r2876(0 to 0));
                                b2894 := ("0" = r2878(0 to 0));
                                b2896 := ("1" = r2880(0 to 0));
                                b2898 := true;
                                b2900 := true;
                                b2902 := true;
                                b2904 := true;
                                b2906 := (b2872 AND (b2890 AND (b2892 AND (b2894 AND (b2896 AND (b2898 AND (b2900 AND (b2902 AND b2904))))))));
                                goto_L2909 := b2906;
                                if (NOT goto_L2909) then
                                  goto_L3057 := (NOT b2906);
                                  null; -- label L3057
                                  -- alt exit (no match)
                                  b3058 := true;
                                  r3060 := r730(0 to 0);
                                  r3062 := r730(1 to 1);
                                  r3064 := r730(2 to 2);
                                  r3066 := r730(3 to 3);
                                  r3068 := r730(4 to 4);
                                  r3070 := r730(5 to 5);
                                  r3072 := r730(6 to 6);
                                  r3074 := r730(7 to 7);
                                  b3076 := ("1" = r3060(0 to 0));
                                  b3078 := ("0" = r3062(0 to 0));
                                  b3080 := ("1" = r3064(0 to 0));
                                  b3082 := ("0" = r3066(0 to 0));
                                  b3084 := true;
                                  b3086 := true;
                                  b3088 := true;
                                  b3090 := true;
                                  b3092 := (b3058 AND (b3076 AND (b3078 AND (b3080 AND (b3082 AND (b3084 AND (b3086 AND (b3088 AND b3090))))))));
                                  goto_L3095 := b3092;
                                  if (NOT goto_L3095) then
                                    goto_L3243 := (NOT b3092);
                                    null; -- label L3243
                                    -- alt exit (no match)
                                    b3244 := true;
                                    r3246 := r730(0 to 0);
                                    r3248 := r730(1 to 1);
                                    r3250 := r730(2 to 2);
                                    r3252 := r730(3 to 3);
                                    r3254 := r730(4 to 4);
                                    r3256 := r730(5 to 5);
                                    r3258 := r730(6 to 6);
                                    r3260 := r730(7 to 7);
                                    b3262 := ("1" = r3246(0 to 0));
                                    b3264 := ("0" = r3248(0 to 0));
                                    b3266 := ("1" = r3250(0 to 0));
                                    b3268 := ("1" = r3252(0 to 0));
                                    b3270 := true;
                                    b3272 := true;
                                    b3274 := true;
                                    b3276 := true;
                                    b3278 := (b3244 AND (b3262 AND (b3264 AND (b3266 AND (b3268 AND (b3270 AND (b3272 AND (b3274 AND b3276))))))));
                                    goto_L3281 := b3278;
                                    if (NOT goto_L3281) then
                                      goto_L3417 := (NOT b3278);
                                      null; -- label L3417
                                      -- alt exit (no match)
                                      b3418 := true;
                                      r3420 := r730(0 to 0);
                                      r3422 := r730(1 to 1);
                                      r3424 := r730(2 to 2);
                                      r3426 := r730(3 to 3);
                                      r3428 := r730(4 to 4);
                                      r3430 := r730(5 to 5);
                                      r3432 := r730(6 to 6);
                                      r3434 := r730(7 to 7);
                                      b3436 := ("1" = r3420(0 to 0));
                                      b3438 := ("1" = r3422(0 to 0));
                                      b3440 := ("0" = r3424(0 to 0));
                                      b3442 := ("0" = r3426(0 to 0));
                                      b3444 := ("0" = r3428(0 to 0));
                                      b3446 := ("0" = r3430(0 to 0));
                                      b3448 := true;
                                      b3450 := true;
                                      b3452 := (b3418 AND (b3436 AND (b3438 AND (b3440 AND (b3442 AND (b3444 AND (b3446 AND (b3448 AND b3450))))))));
                                      goto_L3455 := b3452;
                                      if (NOT goto_L3455) then
                                        goto_L3526 := (NOT b3452);
                                        null; -- label L3526
                                        -- alt exit (no match)
                                        b3527 := true;
                                        r3529 := r730(0 to 0);
                                        r3531 := r730(1 to 1);
                                        r3533 := r730(2 to 2);
                                        r3535 := r730(3 to 3);
                                        r3537 := r730(4 to 4);
                                        r3539 := r730(5 to 5);
                                        r3541 := r730(6 to 6);
                                        r3543 := r730(7 to 7);
                                        b3545 := ("1" = r3529(0 to 0));
                                        b3547 := ("1" = r3531(0 to 0));
                                        b3549 := ("0" = r3533(0 to 0));
                                        b3551 := ("0" = r3535(0 to 0));
                                        b3553 := ("0" = r3537(0 to 0));
                                        b3555 := ("1" = r3539(0 to 0));
                                        b3557 := true;
                                        b3559 := true;
                                        b3561 := (b3527 AND (b3545 AND (b3547 AND (b3549 AND (b3551 AND (b3553 AND (b3555 AND (b3557 AND b3559))))))));
                                        goto_L3564 := b3561;
                                        if (NOT goto_L3564) then
                                          goto_L3637 := (NOT b3561);
                                          null; -- label L3637
                                          -- alt exit (no match)
                                          b3638 := true;
                                          r3640 := r730(0 to 0);
                                          r3642 := r730(1 to 1);
                                          r3644 := r730(2 to 2);
                                          r3646 := r730(3 to 3);
                                          r3648 := r730(4 to 4);
                                          r3650 := r730(5 to 5);
                                          r3652 := r730(6 to 6);
                                          r3654 := r730(7 to 7);
                                          b3656 := ("1" = r3640(0 to 0));
                                          b3658 := ("1" = r3642(0 to 0));
                                          b3660 := ("0" = r3644(0 to 0));
                                          b3662 := ("0" = r3646(0 to 0));
                                          b3664 := ("1" = r3648(0 to 0));
                                          b3666 := ("0" = r3650(0 to 0));
                                          b3668 := true;
                                          b3670 := true;
                                          b3672 := (b3638 AND (b3656 AND (b3658 AND (b3660 AND (b3662 AND (b3664 AND (b3666 AND (b3668 AND b3670))))))));
                                          goto_L3675 := b3672;
                                          if (NOT goto_L3675) then
                                            goto_L3746 := (NOT b3672);
                                            null; -- label L3746
                                            -- alt exit (no match)
                                            b3747 := true;
                                            r3749 := r730(0 to 0);
                                            r3751 := r730(1 to 1);
                                            r3753 := r730(2 to 2);
                                            r3755 := r730(3 to 3);
                                            r3757 := r730(4 to 4);
                                            r3759 := r730(5 to 5);
                                            r3761 := r730(6 to 6);
                                            r3763 := r730(7 to 7);
                                            b3765 := ("1" = r3749(0 to 0));
                                            b3767 := ("1" = r3751(0 to 0));
                                            b3769 := ("0" = r3753(0 to 0));
                                            b3771 := ("0" = r3755(0 to 0));
                                            b3773 := ("1" = r3757(0 to 0));
                                            b3775 := ("1" = r3759(0 to 0));
                                            b3777 := true;
                                            b3779 := true;
                                            b3781 := (b3747 AND (b3765 AND (b3767 AND (b3769 AND (b3771 AND (b3773 AND (b3775 AND (b3777 AND b3779))))))));
                                            goto_L3784 := b3781;
                                            if (NOT goto_L3784) then
                                              goto_L3857 := (NOT b3781);
                                              null; -- label L3857
                                              -- alt exit (no match)
                                              b3858 := true;
                                              r3860 := r730(0 to 0);
                                              r3862 := r730(1 to 1);
                                              r3864 := r730(2 to 2);
                                              r3866 := r730(3 to 3);
                                              r3868 := r730(4 to 4);
                                              r3870 := r730(5 to 5);
                                              r3872 := r730(6 to 6);
                                              r3874 := r730(7 to 7);
                                              b3876 := ("1" = r3860(0 to 0));
                                              b3878 := ("1" = r3862(0 to 0));
                                              b3880 := ("0" = r3864(0 to 0));
                                              b3882 := ("1" = r3866(0 to 0));
                                              b3884 := ("0" = r3868(0 to 0));
                                              b3886 := ("0" = r3870(0 to 0));
                                              b3888 := true;
                                              b3890 := true;
                                              b3892 := (b3858 AND (b3876 AND (b3878 AND (b3880 AND (b3882 AND (b3884 AND (b3886 AND (b3888 AND b3890))))))));
                                              goto_L3895 := b3892;
                                              if (NOT goto_L3895) then
                                                goto_L3952 := (NOT b3892);
                                                null; -- label L3952
                                                -- alt exit (no match)
                                                b3953 := true;
                                                r3955 := r730(0 to 0);
                                                r3957 := r730(1 to 1);
                                                r3959 := r730(2 to 2);
                                                r3961 := r730(3 to 3);
                                                r3963 := r730(4 to 4);
                                                r3965 := r730(5 to 5);
                                                r3967 := r730(6 to 6);
                                                r3969 := r730(7 to 7);
                                                b3971 := ("1" = r3955(0 to 0));
                                                b3973 := ("1" = r3957(0 to 0));
                                                b3975 := ("0" = r3959(0 to 0));
                                                b3977 := ("1" = r3961(0 to 0));
                                                b3979 := ("0" = r3963(0 to 0));
                                                b3981 := ("1" = r3965(0 to 0));
                                                b3983 := ("0" = r3967(0 to 0));
                                                b3985 := true;
                                                b3987 := (b3953 AND (b3971 AND (b3973 AND (b3975 AND (b3977 AND (b3979 AND (b3981 AND (b3983 AND b3985))))))));
                                                goto_L3990 := b3987;
                                                if (NOT goto_L3990) then
                                                  goto_L4013 := (NOT b3987);
                                                  null; -- label L4013
                                                  -- alt exit (no match)
                                                  b4014 := true;
                                                  r4016 := r730(0 to 0);
                                                  r4018 := r730(1 to 1);
                                                  r4020 := r730(2 to 2);
                                                  r4022 := r730(3 to 3);
                                                  r4024 := r730(4 to 4);
                                                  r4026 := r730(5 to 5);
                                                  r4028 := r730(6 to 6);
                                                  r4030 := r730(7 to 7);
                                                  b4032 := ("1" = r4016(0 to 0));
                                                  b4034 := ("1" = r4018(0 to 0));
                                                  b4036 := ("0" = r4020(0 to 0));
                                                  b4038 := ("1" = r4022(0 to 0));
                                                  b4040 := ("0" = r4024(0 to 0));
                                                  b4042 := ("1" = r4026(0 to 0));
                                                  b4044 := ("1" = r4028(0 to 0));
                                                  b4046 := ("0" = r4030(0 to 0));
                                                  b4048 := (b4014 AND (b4032 AND (b4034 AND (b4036 AND (b4038 AND (b4040 AND (b4042 AND (b4044 AND b4046))))))));
                                                  goto_L4051 := b4048;
                                                  if (NOT goto_L4051) then
                                                    goto_L4100 := (NOT b4048);
                                                    null; -- label L4100
                                                    -- alt exit (no match)
                                                    b4101 := true;
                                                    r4103 := r730(0 to 0);
                                                    r4105 := r730(1 to 1);
                                                    r4107 := r730(2 to 2);
                                                    r4109 := r730(3 to 3);
                                                    r4111 := r730(4 to 4);
                                                    r4113 := r730(5 to 5);
                                                    r4115 := r730(6 to 6);
                                                    r4117 := r730(7 to 7);
                                                    b4119 := ("1" = r4103(0 to 0));
                                                    b4121 := ("1" = r4105(0 to 0));
                                                    b4123 := ("0" = r4107(0 to 0));
                                                    b4125 := ("1" = r4109(0 to 0));
                                                    b4127 := ("0" = r4111(0 to 0));
                                                    b4129 := ("1" = r4113(0 to 0));
                                                    b4131 := ("1" = r4115(0 to 0));
                                                    b4133 := ("1" = r4117(0 to 0));
                                                    b4135 := (b4101 AND (b4119 AND (b4121 AND (b4123 AND (b4125 AND (b4127 AND (b4129 AND (b4131 AND b4133))))))));
                                                    goto_L4138 := b4135;
                                                    if (NOT goto_L4138) then
                                                      goto_L4294 := (NOT b4135);
                                                      null; -- label L4294
                                                      -- alt exit (no match)
                                                      b4295 := true;
                                                      r4297 := r730(0 to 0);
                                                      r4299 := r730(1 to 1);
                                                      r4301 := r730(2 to 2);
                                                      r4303 := r730(3 to 3);
                                                      r4305 := r730(4 to 4);
                                                      r4307 := r730(5 to 5);
                                                      r4309 := r730(6 to 6);
                                                      r4311 := r730(7 to 7);
                                                      b4313 := ("1" = r4297(0 to 0));
                                                      b4315 := ("1" = r4299(0 to 0));
                                                      b4317 := ("0" = r4301(0 to 0));
                                                      b4319 := ("1" = r4303(0 to 0));
                                                      b4321 := ("1" = r4305(0 to 0));
                                                      b4323 := ("0" = r4307(0 to 0));
                                                      b4325 := true;
                                                      b4327 := true;
                                                      b4329 := (b4295 AND (b4313 AND (b4315 AND (b4317 AND (b4319 AND (b4321 AND (b4323 AND (b4325 AND b4327))))))));
                                                      goto_L4332 := b4329;
                                                      if (NOT goto_L4332) then
                                                        goto_L4431 := (NOT b4329);
                                                        null; -- label L4431
                                                        -- alt exit (no match)
                                                        b4432 := true;
                                                        r4434 := r730(0 to 0);
                                                        r4436 := r730(1 to 1);
                                                        r4438 := r730(2 to 2);
                                                        r4440 := r730(3 to 3);
                                                        r4442 := r730(4 to 4);
                                                        r4444 := r730(5 to 5);
                                                        r4446 := r730(6 to 6);
                                                        r4448 := r730(7 to 7);
                                                        b4450 := ("1" = r4434(0 to 0));
                                                        b4452 := ("1" = r4436(0 to 0));
                                                        b4454 := ("0" = r4438(0 to 0));
                                                        b4456 := ("1" = r4440(0 to 0));
                                                        b4458 := ("1" = r4442(0 to 0));
                                                        b4460 := ("1" = r4444(0 to 0));
                                                        b4462 := true;
                                                        b4464 := true;
                                                        b4466 := (b4432 AND (b4450 AND (b4452 AND (b4454 AND (b4456 AND (b4458 AND (b4460 AND (b4462 AND b4464))))))));
                                                        goto_L4469 := b4466;
                                                        if (NOT goto_L4469) then
                                                          goto_L4530 := (NOT b4466);
                                                          null; -- label L4530
                                                          -- alt exit (no match)
                                                          b4531 := true;
                                                          r4533 := r730(0 to 0);
                                                          r4535 := r730(1 to 1);
                                                          r4537 := r730(2 to 2);
                                                          r4539 := r730(3 to 3);
                                                          r4541 := r730(4 to 4);
                                                          r4543 := r730(5 to 5);
                                                          r4545 := r730(6 to 6);
                                                          r4547 := r730(7 to 7);
                                                          b4549 := ("1" = r4533(0 to 0));
                                                          b4551 := ("1" = r4535(0 to 0));
                                                          b4553 := ("1" = r4537(0 to 0));
                                                          b4555 := ("0" = r4539(0 to 0));
                                                          b4557 := ("0" = r4541(0 to 0));
                                                          b4559 := ("0" = r4543(0 to 0));
                                                          b4561 := true;
                                                          b4563 := true;
                                                          b4565 := (b4531 AND (b4549 AND (b4551 AND (b4553 AND (b4555 AND (b4557 AND (b4559 AND (b4561 AND b4563))))))));
                                                          goto_L4568 := b4565;
                                                          if (NOT goto_L4568) then
                                                            goto_L4712 := (NOT b4565);
                                                            null; -- label L4712
                                                            -- alt exit (no match)
                                                            b4713 := true;
                                                            r4715 := r730(0 to 0);
                                                            r4717 := r730(1 to 1);
                                                            r4719 := r730(2 to 2);
                                                            r4721 := r730(3 to 3);
                                                            r4723 := r730(4 to 4);
                                                            r4725 := r730(5 to 5);
                                                            r4727 := r730(6 to 6);
                                                            r4729 := r730(7 to 7);
                                                            b4731 := ("1" = r4715(0 to 0));
                                                            b4733 := ("1" = r4717(0 to 0));
                                                            b4735 := ("1" = r4719(0 to 0));
                                                            b4737 := ("0" = r4721(0 to 0));
                                                            b4739 := ("0" = r4723(0 to 0));
                                                            b4741 := ("1" = r4725(0 to 0));
                                                            b4743 := true;
                                                            b4745 := true;
                                                            b4747 := (b4713 AND (b4731 AND (b4733 AND (b4735 AND (b4737 AND (b4739 AND (b4741 AND (b4743 AND b4745))))))));
                                                            goto_L4750 := b4747;
                                                            if (NOT goto_L4750) then
                                                              goto_L4894 := (NOT b4747);
                                                              null; -- label L4894
                                                              -- alt exit (no match)
                                                              b4895 := true;
                                                              r4897 := r730(0 to 0);
                                                              r4899 := r730(1 to 1);
                                                              r4901 := r730(2 to 2);
                                                              r4903 := r730(3 to 3);
                                                              r4905 := r730(4 to 4);
                                                              r4907 := r730(5 to 5);
                                                              r4909 := r730(6 to 6);
                                                              r4911 := r730(7 to 7);
                                                              b4913 := ("1" = r4897(0 to 0));
                                                              b4915 := ("1" = r4899(0 to 0));
                                                              b4917 := ("1" = r4901(0 to 0));
                                                              b4919 := ("0" = r4903(0 to 0));
                                                              b4921 := ("1" = r4905(0 to 0));
                                                              b4923 := true;
                                                              b4925 := true;
                                                              b4927 := true;
                                                              b4929 := (b4895 AND (b4913 AND (b4915 AND (b4917 AND (b4919 AND (b4921 AND (b4923 AND (b4925 AND b4927))))))));
                                                              goto_L4931 := b4929;
                                                              if (NOT goto_L4931) then
                                                                goto_L5138 := (NOT b4929);
                                                                null; -- label L5138
                                                                -- alt exit (no match)
                                                                b5139 := true;
                                                                r5141 := r730(0 to 0);
                                                                r5143 := r730(1 to 1);
                                                                r5145 := r730(2 to 2);
                                                                r5147 := r730(3 to 3);
                                                                r5149 := r730(4 to 4);
                                                                r5151 := r730(5 to 5);
                                                                r5153 := r730(6 to 6);
                                                                r5155 := r730(7 to 7);
                                                                b5157 := ("1" = r5141(0 to 0));
                                                                b5159 := ("1" = r5143(0 to 0));
                                                                b5161 := ("1" = r5145(0 to 0));
                                                                b5163 := ("1" = r5147(0 to 0));
                                                                b5165 := true;
                                                                b5167 := true;
                                                                b5169 := true;
                                                                b5171 := true;
                                                                b5173 := (b5139 AND (b5157 AND (b5159 AND (b5161 AND (b5163 AND (b5165 AND (b5167 AND (b5169 AND b5171))))))));
                                                                goto_L5176 := b5173;
                                                                if (NOT goto_L5176) then
                                                                  goto_L5392 := (NOT b5173);
                                                                  null; -- label L5392
                                                                  -- alt exit (no match)
                                                                  b5393 := true;
                                                                  r5395 := statevar0;
                                                                  -- got s@MN in r5395
                                                                  r5398 := "0";
                                                                  r5400 := rewire_setCFlag_5(r5395,r5398);
                                                                  statevar0 := r5400;
                                                                  r5403 := statevar0;
                                                                  -- got s@MP in r5403
                                                                  r5406 := "0";
                                                                  r5408 := rewire_setZFlag_48(r5403,r5406);
                                                                  statevar0 := r5408;
                                                                  r5411 := statevar0;
                                                                  -- got s@MR in r5411
                                                                  r5414 := rewire_initOutputs_127;
                                                                  r5416 := rewire_setOutputs_91(r5411,r5414);
                                                                  statevar0 := r5416;
                                                                  r5419 := statevar0;
                                                                  -- got s@MT in r5419
                                                                  r5422 := rewire_outputs_144(r5419);
                                                                  -- got o@MU in r5422
                                                                  nextout := r5422;
                                                                  state := STATE5427;
                                                                  goto_L5439 := true;
                                                                end if;
                                                                goto_L5439 := goto_L5439;
                                                                if (NOT goto_L5439) then
                                                                  null; -- label L5176
                                                                  r5175 := statevar0;
                                                                  -- got b0@M4 in r5153
                                                                  -- got b1@M5 in r5155
                                                                  r5179 := rewire_mkReg_883(r5153,r5155);
                                                                  b5183 := ("00" = r5179(0 to 1));
                                                                  goto_L5185 := b5183;
                                                                  if (NOT goto_L5185) then
                                                                    goto_L5189 := (NOT b5183);
                                                                    null; -- label L5189
                                                                    -- alt exit (no match)
                                                                    b5190 := ("01" = r5179(0 to 1));
                                                                    goto_L5192 := b5190;
                                                                    if (NOT goto_L5192) then
                                                                      goto_L5196 := (NOT b5190);
                                                                      null; -- label L5196
                                                                      -- alt exit (no match)
                                                                      b5197 := ("10" = r5179(0 to 1));
                                                                      goto_L5199 := b5197;
                                                                      if (NOT goto_L5199) then
                                                                        goto_L5203 := (NOT b5197);
                                                                        null; -- label L5203
                                                                        -- alt exit (no match)
                                                                        -- final pat
                                                                        -- got s@M6 in r5175
                                                                        r5206 := rewire_r3_1046(r5175);
                                                                        r5181 := r5206;
                                                                        goto_L5182 := true;
                                                                      end if;
                                                                      goto_L5182 := goto_L5182;
                                                                      if (NOT goto_L5182) then
                                                                        null; -- label L5199
                                                                        -- got s@M6 in r5175
                                                                        r5200 := rewire_r2_1008(r5175);
                                                                        r5181 := r5200;
                                                                        goto_L5182 := true;
                                                                      end if;
                                                                      goto_L5182 := goto_L5182;
                                                                    end if;
                                                                    goto_L5182 := goto_L5182;
                                                                    if (NOT goto_L5182) then
                                                                      null; -- label L5192
                                                                      -- got s@M6 in r5175
                                                                      r5193 := rewire_r1_969(r5175);
                                                                      r5181 := r5193;
                                                                      goto_L5182 := true;
                                                                    end if;
                                                                    goto_L5182 := goto_L5182;
                                                                  end if;
                                                                  goto_L5182 := goto_L5182;
                                                                  if (NOT goto_L5182) then
                                                                    null; -- label L5185
                                                                    -- got s@M6 in r5175
                                                                    r5186 := rewire_r0_930(r5175);
                                                                    r5181 := r5186;
                                                                    goto_L5182 := true;
                                                                  end if;
                                                                  goto_L5182 := goto_L5182;
                                                                  null; -- label L5182
                                                                  -- end case
                                                                  null;
                                                                  -- got d@M3 in r5151
                                                                  -- got l@M2 in r5149
                                                                  r5212 := (r5151 & r5149);
                                                                  b5215 := true;
                                                                  r5217 := r5212(0 to 0);
                                                                  r5219 := r5212(1 to 1);
                                                                  b5221 := ("0" = r5217(0 to 0));
                                                                  b5223 := ("0" = r5219(0 to 0));
                                                                  b5225 := (b5215 AND (b5221 AND b5223));
                                                                  goto_L5227 := b5225;
                                                                  if (NOT goto_L5227) then
                                                                    goto_L5234 := (NOT b5225);
                                                                    null; -- label L5234
                                                                    -- alt exit (no match)
                                                                    b5235 := true;
                                                                    r5237 := r5212(0 to 0);
                                                                    r5239 := r5212(1 to 1);
                                                                    b5241 := ("0" = r5237(0 to 0));
                                                                    b5243 := ("1" = r5239(0 to 0));
                                                                    b5245 := (b5235 AND (b5241 AND b5243));
                                                                    goto_L5247 := b5245;
                                                                    if (NOT goto_L5247) then
                                                                      goto_L5253 := (NOT b5245);
                                                                      null; -- label L5253
                                                                      -- alt exit (no match)
                                                                      b5254 := true;
                                                                      r5256 := r5212(0 to 0);
                                                                      r5258 := r5212(1 to 1);
                                                                      b5260 := ("1" = r5256(0 to 0));
                                                                      b5262 := ("0" = r5258(0 to 0));
                                                                      b5264 := (b5254 AND (b5260 AND b5262));
                                                                      goto_L5266 := b5264;
                                                                      if (NOT goto_L5266) then
                                                                        goto_L5273 := (NOT b5264);
                                                                        null; -- label L5273
                                                                        -- alt exit (no match)
                                                                        -- final pat
                                                                        r5275 := r5212(0 to 0);
                                                                        r5277 := r5212(1 to 1);
                                                                        -- final pat
                                                                        -- final pat
                                                                        -- got v@M7 in r5181
                                                                        r5282 := "0";
                                                                        r5284 := shrCW8(r5181,r5282);
                                                                        r5214 := r5284;
                                                                        goto_L5287 := true;
                                                                      end if;
                                                                      goto_L5287 := goto_L5287;
                                                                      if (NOT goto_L5287) then
                                                                        null; -- label L5266
                                                                        -- got v@M7 in r5181
                                                                        -- got v@M7 in r5181
                                                                        r5268 := lsbW8(r5181);
                                                                        r5270 := shrCW8(r5181,r5268);
                                                                        r5214 := r5270;
                                                                        goto_L5287 := true;
                                                                      end if;
                                                                      goto_L5287 := goto_L5287;
                                                                    end if;
                                                                    goto_L5287 := goto_L5287;
                                                                    if (NOT goto_L5287) then
                                                                      null; -- label L5247
                                                                      -- got v@M7 in r5181
                                                                      r5248 := "0";
                                                                      r5250 := shlCW8(r5181,r5248);
                                                                      r5214 := r5250;
                                                                      goto_L5287 := true;
                                                                    end if;
                                                                    goto_L5287 := goto_L5287;
                                                                  end if;
                                                                  goto_L5287 := goto_L5287;
                                                                  if (NOT goto_L5287) then
                                                                    null; -- label L5227
                                                                    -- got v@M7 in r5181
                                                                    -- got v@M7 in r5181
                                                                    r5229 := msbW8(r5181);
                                                                    r5231 := shlCW8(r5181,r5229);
                                                                    r5214 := r5231;
                                                                    goto_L5287 := true;
                                                                  end if;
                                                                  goto_L5287 := goto_L5287;
                                                                  null; -- label L5287
                                                                  -- end case
                                                                  -- got p@M8 in r5214
                                                                  -- final pat
                                                                  r5291 := r5214(0 to 0);
                                                                  r5293 := r5214(1 to 8);
                                                                  b5295 := true;
                                                                  b5297 := true;
                                                                  -- got x@M9 in r5291
                                                                  r5289 := r5291;
                                                                  -- end case
                                                                  -- got p@M8 in r5214
                                                                  -- final pat
                                                                  r5305 := r5214(0 to 0);
                                                                  r5307 := r5214(1 to 8);
                                                                  b5309 := true;
                                                                  b5311 := true;
                                                                  -- got x@MB in r5307
                                                                  r5303 := r5307;
                                                                  -- end case
                                                                  r5316 := statevar0;
                                                                  -- got b0@M4 in r5153
                                                                  -- got b1@M5 in r5155
                                                                  r5320 := rewire_mkReg_883(r5153,r5155);
                                                                  b5323 := ("00" = r5320(0 to 1));
                                                                  goto_L5325 := b5323;
                                                                  if (NOT goto_L5325) then
                                                                    goto_L5331 := (NOT b5323);
                                                                    null; -- label L5331
                                                                    -- alt exit (no match)
                                                                    b5332 := ("01" = r5320(0 to 1));
                                                                    goto_L5334 := b5332;
                                                                    if (NOT goto_L5334) then
                                                                      goto_L5340 := (NOT b5332);
                                                                      null; -- label L5340
                                                                      -- alt exit (no match)
                                                                      b5341 := ("10" = r5320(0 to 1));
                                                                      goto_L5343 := b5341;
                                                                      if (NOT goto_L5343) then
                                                                        goto_L5349 := (NOT b5341);
                                                                        null; -- label L5349
                                                                        -- alt exit (no match)
                                                                        -- final pat
                                                                        -- got s@MD in r5316
                                                                        -- got v'@MC in r5303
                                                                        r5353 := rewire_setR3_1349(r5316,r5303);
                                                                        statevar0 := r5353;
                                                                        null;
                                                                        goto_L5322 := true;
                                                                      end if;
                                                                      goto_L5322 := goto_L5322;
                                                                      if (NOT goto_L5322) then
                                                                        null; -- label L5343
                                                                        -- got s@MD in r5316
                                                                        -- got v'@MC in r5303
                                                                        r5345 := rewire_setR2_1306(r5316,r5303);
                                                                        statevar0 := r5345;
                                                                        null;
                                                                        goto_L5322 := true;
                                                                      end if;
                                                                      goto_L5322 := goto_L5322;
                                                                    end if;
                                                                    goto_L5322 := goto_L5322;
                                                                    if (NOT goto_L5322) then
                                                                      null; -- label L5334
                                                                      -- got s@MD in r5316
                                                                      -- got v'@MC in r5303
                                                                      r5336 := rewire_setR1_1262(r5316,r5303);
                                                                      statevar0 := r5336;
                                                                      null;
                                                                      goto_L5322 := true;
                                                                    end if;
                                                                    goto_L5322 := goto_L5322;
                                                                  end if;
                                                                  goto_L5322 := goto_L5322;
                                                                  if (NOT goto_L5322) then
                                                                    null; -- label L5325
                                                                    -- got s@MD in r5316
                                                                    -- got v'@MC in r5303
                                                                    r5327 := rewire_setR0_1218(r5316,r5303);
                                                                    statevar0 := r5327;
                                                                    null;
                                                                    goto_L5322 := true;
                                                                  end if;
                                                                  goto_L5322 := goto_L5322;
                                                                  null; -- label L5322
                                                                  -- end case
                                                                  r5357 := statevar0;
                                                                  -- got s@MF in r5357
                                                                  -- got cout@MA in r5289
                                                                  r5361 := rewire_setCFlag_5(r5357,r5289);
                                                                  statevar0 := r5361;
                                                                  r5364 := statevar0;
                                                                  -- got s@MH in r5364
                                                                  -- got v'@MC in r5303
                                                                  r5368 := zeroW8;
                                                                  r5370 := eqW8(r5303,r5368);
                                                                  r5372 := rewire_setZFlag_48(r5364,r5370);
                                                                  statevar0 := r5372;
                                                                  r5375 := statevar0;
                                                                  -- got s@MJ in r5375
                                                                  r5378 := rewire_outputs_144(r5375);
                                                                  -- got o@MK in r5378
                                                                  nextout := r5378;
                                                                  state := STATE5383;
                                                                  goto_L5439 := true;
                                                                end if;
                                                                goto_L5439 := goto_L5439;
                                                              end if;
                                                              goto_L5439 := goto_L5439;
                                                              if (NOT goto_L5439) then
                                                                null; -- label L4931
                                                                -- got d@LF in r4907
                                                                b4933 := ("0" = r4907(0 to 0));
                                                                goto_L4936 := b4933;
                                                                if (NOT goto_L4936) then
                                                                  goto_L5035 := (NOT b4933);
                                                                  null; -- label L5035
                                                                  -- alt exit (no match)
                                                                  -- final pat
                                                                  r5037 := statevar0;
                                                                  -- got b0@LG in r4909
                                                                  -- got b1@LH in r4911
                                                                  r5041 := rewire_mkReg_883(r4909,r4911);
                                                                  b5045 := ("00" = r5041(0 to 1));
                                                                  goto_L5047 := b5045;
                                                                  if (NOT goto_L5047) then
                                                                    goto_L5051 := (NOT b5045);
                                                                    null; -- label L5051
                                                                    -- alt exit (no match)
                                                                    b5052 := ("01" = r5041(0 to 1));
                                                                    goto_L5054 := b5052;
                                                                    if (NOT goto_L5054) then
                                                                      goto_L5058 := (NOT b5052);
                                                                      null; -- label L5058
                                                                      -- alt exit (no match)
                                                                      b5059 := ("10" = r5041(0 to 1));
                                                                      goto_L5061 := b5059;
                                                                      if (NOT goto_L5061) then
                                                                        goto_L5065 := (NOT b5059);
                                                                        null; -- label L5065
                                                                        -- alt exit (no match)
                                                                        -- final pat
                                                                        -- got s@LQ in r5037
                                                                        r5068 := rewire_r3_1046(r5037);
                                                                        r5043 := r5068;
                                                                        goto_L5044 := true;
                                                                      end if;
                                                                      goto_L5044 := goto_L5044;
                                                                      if (NOT goto_L5044) then
                                                                        null; -- label L5061
                                                                        -- got s@LQ in r5037
                                                                        r5062 := rewire_r2_1008(r5037);
                                                                        r5043 := r5062;
                                                                        goto_L5044 := true;
                                                                      end if;
                                                                      goto_L5044 := goto_L5044;
                                                                    end if;
                                                                    goto_L5044 := goto_L5044;
                                                                    if (NOT goto_L5044) then
                                                                      null; -- label L5054
                                                                      -- got s@LQ in r5037
                                                                      r5055 := rewire_r1_969(r5037);
                                                                      r5043 := r5055;
                                                                      goto_L5044 := true;
                                                                    end if;
                                                                    goto_L5044 := goto_L5044;
                                                                  end if;
                                                                  goto_L5044 := goto_L5044;
                                                                  if (NOT goto_L5044) then
                                                                    null; -- label L5047
                                                                    -- got s@LQ in r5037
                                                                    r5048 := rewire_r0_930(r5037);
                                                                    r5043 := r5048;
                                                                    goto_L5044 := true;
                                                                  end if;
                                                                  goto_L5044 := goto_L5044;
                                                                  null; -- label L5044
                                                                  -- end case
                                                                  r5071 := statevar0;
                                                                  -- got b0@LG in r4909
                                                                  -- got b1@LH in r4911
                                                                  r5075 := rewire_mkReg_883(r4909,r4911);
                                                                  b5078 := ("00" = r5075(0 to 1));
                                                                  goto_L5080 := b5078;
                                                                  if (NOT goto_L5080) then
                                                                    goto_L5088 := (NOT b5078);
                                                                    null; -- label L5088
                                                                    -- alt exit (no match)
                                                                    b5089 := ("01" = r5075(0 to 1));
                                                                    goto_L5091 := b5089;
                                                                    if (NOT goto_L5091) then
                                                                      goto_L5099 := (NOT b5089);
                                                                      null; -- label L5099
                                                                      -- alt exit (no match)
                                                                      b5100 := ("10" = r5075(0 to 1));
                                                                      goto_L5102 := b5100;
                                                                      if (NOT goto_L5102) then
                                                                        goto_L5110 := (NOT b5100);
                                                                        null; -- label L5110
                                                                        -- alt exit (no match)
                                                                        -- final pat
                                                                        -- got s@LS in r5071
                                                                        -- got v@LR in r5043
                                                                        r5114 := rorW8(r5043);
                                                                        r5116 := rewire_setR3_1349(r5071,r5114);
                                                                        statevar0 := r5116;
                                                                        null;
                                                                        goto_L5077 := true;
                                                                      end if;
                                                                      goto_L5077 := goto_L5077;
                                                                      if (NOT goto_L5077) then
                                                                        null; -- label L5102
                                                                        -- got s@LS in r5071
                                                                        -- got v@LR in r5043
                                                                        r5104 := rorW8(r5043);
                                                                        r5106 := rewire_setR2_1306(r5071,r5104);
                                                                        statevar0 := r5106;
                                                                        null;
                                                                        goto_L5077 := true;
                                                                      end if;
                                                                      goto_L5077 := goto_L5077;
                                                                    end if;
                                                                    goto_L5077 := goto_L5077;
                                                                    if (NOT goto_L5077) then
                                                                      null; -- label L5091
                                                                      -- got s@LS in r5071
                                                                      -- got v@LR in r5043
                                                                      r5093 := rorW8(r5043);
                                                                      r5095 := rewire_setR1_1262(r5071,r5093);
                                                                      statevar0 := r5095;
                                                                      null;
                                                                      goto_L5077 := true;
                                                                    end if;
                                                                    goto_L5077 := goto_L5077;
                                                                  end if;
                                                                  goto_L5077 := goto_L5077;
                                                                  if (NOT goto_L5077) then
                                                                    null; -- label L5080
                                                                    -- got s@LS in r5071
                                                                    -- got v@LR in r5043
                                                                    r5082 := rorW8(r5043);
                                                                    r5084 := rewire_setR0_1218(r5071,r5082);
                                                                    statevar0 := r5084;
                                                                    null;
                                                                    goto_L5077 := true;
                                                                  end if;
                                                                  goto_L5077 := goto_L5077;
                                                                  null; -- label L5077
                                                                  -- end case
                                                                  r5120 := statevar0;
                                                                  -- got s@LU in r5120
                                                                  r5123 := rewire_outputs_144(r5120);
                                                                  -- got o@LV in r5123
                                                                  nextout := r5123;
                                                                  state := STATE5128;
                                                                  goto_L5439 := true;
                                                                end if;
                                                                goto_L5439 := goto_L5439;
                                                                if (NOT goto_L5439) then
                                                                  null; -- label L4936
                                                                  r4935 := statevar0;
                                                                  -- got b0@LG in r4909
                                                                  -- got b1@LH in r4911
                                                                  r4939 := rewire_mkReg_883(r4909,r4911);
                                                                  b4943 := ("00" = r4939(0 to 1));
                                                                  goto_L4945 := b4943;
                                                                  if (NOT goto_L4945) then
                                                                    goto_L4949 := (NOT b4943);
                                                                    null; -- label L4949
                                                                    -- alt exit (no match)
                                                                    b4950 := ("01" = r4939(0 to 1));
                                                                    goto_L4952 := b4950;
                                                                    if (NOT goto_L4952) then
                                                                      goto_L4956 := (NOT b4950);
                                                                      null; -- label L4956
                                                                      -- alt exit (no match)
                                                                      b4957 := ("10" = r4939(0 to 1));
                                                                      goto_L4959 := b4957;
                                                                      if (NOT goto_L4959) then
                                                                        goto_L4963 := (NOT b4957);
                                                                        null; -- label L4963
                                                                        -- alt exit (no match)
                                                                        -- final pat
                                                                        -- got s@LI in r4935
                                                                        r4966 := rewire_r3_1046(r4935);
                                                                        r4941 := r4966;
                                                                        goto_L4942 := true;
                                                                      end if;
                                                                      goto_L4942 := goto_L4942;
                                                                      if (NOT goto_L4942) then
                                                                        null; -- label L4959
                                                                        -- got s@LI in r4935
                                                                        r4960 := rewire_r2_1008(r4935);
                                                                        r4941 := r4960;
                                                                        goto_L4942 := true;
                                                                      end if;
                                                                      goto_L4942 := goto_L4942;
                                                                    end if;
                                                                    goto_L4942 := goto_L4942;
                                                                    if (NOT goto_L4942) then
                                                                      null; -- label L4952
                                                                      -- got s@LI in r4935
                                                                      r4953 := rewire_r1_969(r4935);
                                                                      r4941 := r4953;
                                                                      goto_L4942 := true;
                                                                    end if;
                                                                    goto_L4942 := goto_L4942;
                                                                  end if;
                                                                  goto_L4942 := goto_L4942;
                                                                  if (NOT goto_L4942) then
                                                                    null; -- label L4945
                                                                    -- got s@LI in r4935
                                                                    r4946 := rewire_r0_930(r4935);
                                                                    r4941 := r4946;
                                                                    goto_L4942 := true;
                                                                  end if;
                                                                  goto_L4942 := goto_L4942;
                                                                  null; -- label L4942
                                                                  -- end case
                                                                  r4969 := statevar0;
                                                                  -- got b0@LG in r4909
                                                                  -- got b1@LH in r4911
                                                                  r4973 := rewire_mkReg_883(r4909,r4911);
                                                                  b4976 := ("00" = r4973(0 to 1));
                                                                  goto_L4978 := b4976;
                                                                  if (NOT goto_L4978) then
                                                                    goto_L4986 := (NOT b4976);
                                                                    null; -- label L4986
                                                                    -- alt exit (no match)
                                                                    b4987 := ("01" = r4973(0 to 1));
                                                                    goto_L4989 := b4987;
                                                                    if (NOT goto_L4989) then
                                                                      goto_L4997 := (NOT b4987);
                                                                      null; -- label L4997
                                                                      -- alt exit (no match)
                                                                      b4998 := ("10" = r4973(0 to 1));
                                                                      goto_L5000 := b4998;
                                                                      if (NOT goto_L5000) then
                                                                        goto_L5008 := (NOT b4998);
                                                                        null; -- label L5008
                                                                        -- alt exit (no match)
                                                                        -- final pat
                                                                        -- got s@LK in r4969
                                                                        -- got v@LJ in r4941
                                                                        r5012 := rolW8(r4941);
                                                                        r5014 := rewire_setR3_1349(r4969,r5012);
                                                                        statevar0 := r5014;
                                                                        null;
                                                                        goto_L4975 := true;
                                                                      end if;
                                                                      goto_L4975 := goto_L4975;
                                                                      if (NOT goto_L4975) then
                                                                        null; -- label L5000
                                                                        -- got s@LK in r4969
                                                                        -- got v@LJ in r4941
                                                                        r5002 := rolW8(r4941);
                                                                        r5004 := rewire_setR2_1306(r4969,r5002);
                                                                        statevar0 := r5004;
                                                                        null;
                                                                        goto_L4975 := true;
                                                                      end if;
                                                                      goto_L4975 := goto_L4975;
                                                                    end if;
                                                                    goto_L4975 := goto_L4975;
                                                                    if (NOT goto_L4975) then
                                                                      null; -- label L4989
                                                                      -- got s@LK in r4969
                                                                      -- got v@LJ in r4941
                                                                      r4991 := rolW8(r4941);
                                                                      r4993 := rewire_setR1_1262(r4969,r4991);
                                                                      statevar0 := r4993;
                                                                      null;
                                                                      goto_L4975 := true;
                                                                    end if;
                                                                    goto_L4975 := goto_L4975;
                                                                  end if;
                                                                  goto_L4975 := goto_L4975;
                                                                  if (NOT goto_L4975) then
                                                                    null; -- label L4978
                                                                    -- got s@LK in r4969
                                                                    -- got v@LJ in r4941
                                                                    r4980 := rolW8(r4941);
                                                                    r4982 := rewire_setR0_1218(r4969,r4980);
                                                                    statevar0 := r4982;
                                                                    null;
                                                                    goto_L4975 := true;
                                                                  end if;
                                                                  goto_L4975 := goto_L4975;
                                                                  null; -- label L4975
                                                                  -- end case
                                                                  r5018 := statevar0;
                                                                  -- got s@LM in r5018
                                                                  r5021 := rewire_outputs_144(r5018);
                                                                  -- got o@LN in r5021
                                                                  nextout := r5021;
                                                                  state := STATE5026;
                                                                  goto_L5439 := true;
                                                                end if;
                                                                goto_L5439 := goto_L5439;
                                                              end if;
                                                              goto_L5439 := goto_L5439;
                                                            end if;
                                                            goto_L5439 := goto_L5439;
                                                            if (NOT goto_L5439) then
                                                              null; -- label L4750
                                                              r4749 := statevar0;
                                                              -- got b0@KS in r4727
                                                              -- got b1@KT in r4729
                                                              r4753 := rewire_mkReg_883(r4727,r4729);
                                                              b4757 := ("00" = r4753(0 to 1));
                                                              goto_L4759 := b4757;
                                                              if (NOT goto_L4759) then
                                                                goto_L4763 := (NOT b4757);
                                                                null; -- label L4763
                                                                -- alt exit (no match)
                                                                b4764 := ("01" = r4753(0 to 1));
                                                                goto_L4766 := b4764;
                                                                if (NOT goto_L4766) then
                                                                  goto_L4770 := (NOT b4764);
                                                                  null; -- label L4770
                                                                  -- alt exit (no match)
                                                                  b4771 := ("10" = r4753(0 to 1));
                                                                  goto_L4773 := b4771;
                                                                  if (NOT goto_L4773) then
                                                                    goto_L4777 := (NOT b4771);
                                                                    null; -- label L4777
                                                                    -- alt exit (no match)
                                                                    -- final pat
                                                                    -- got s@KU in r4749
                                                                    r4780 := rewire_r3_1046(r4749);
                                                                    r4755 := r4780;
                                                                    goto_L4756 := true;
                                                                  end if;
                                                                  goto_L4756 := goto_L4756;
                                                                  if (NOT goto_L4756) then
                                                                    null; -- label L4773
                                                                    -- got s@KU in r4749
                                                                    r4774 := rewire_r2_1008(r4749);
                                                                    r4755 := r4774;
                                                                    goto_L4756 := true;
                                                                  end if;
                                                                  goto_L4756 := goto_L4756;
                                                                end if;
                                                                goto_L4756 := goto_L4756;
                                                                if (NOT goto_L4756) then
                                                                  null; -- label L4766
                                                                  -- got s@KU in r4749
                                                                  r4767 := rewire_r1_969(r4749);
                                                                  r4755 := r4767;
                                                                  goto_L4756 := true;
                                                                end if;
                                                                goto_L4756 := goto_L4756;
                                                              end if;
                                                              goto_L4756 := goto_L4756;
                                                              if (NOT goto_L4756) then
                                                                null; -- label L4759
                                                                -- got s@KU in r4749
                                                                r4760 := rewire_r0_930(r4749);
                                                                r4755 := r4760;
                                                                goto_L4756 := true;
                                                              end if;
                                                              goto_L4756 := goto_L4756;
                                                              null; -- label L4756
                                                              -- end case
                                                              -- got v@KV in r4755
                                                              r4784 := oneW8;
                                                              r4786 := "0";
                                                              r4788 := minusCW8(r4755,r4784,r4786);
                                                              -- got p@L0 in r4788
                                                              -- final pat
                                                              r4793 := r4788(0 to 0);
                                                              r4795 := r4788(1 to 8);
                                                              b4797 := true;
                                                              b4799 := true;
                                                              -- got x@L1 in r4793
                                                              r4791 := r4793;
                                                              -- end case
                                                              -- got p@L0 in r4788
                                                              -- final pat
                                                              r4807 := r4788(0 to 0);
                                                              r4809 := r4788(1 to 8);
                                                              b4811 := true;
                                                              b4813 := true;
                                                              -- got x@L3 in r4809
                                                              r4805 := r4809;
                                                              -- end case
                                                              r4818 := statevar0;
                                                              -- got b0@KS in r4727
                                                              -- got b1@KT in r4729
                                                              r4822 := rewire_mkReg_883(r4727,r4729);
                                                              b4825 := ("00" = r4822(0 to 1));
                                                              goto_L4827 := b4825;
                                                              if (NOT goto_L4827) then
                                                                goto_L4833 := (NOT b4825);
                                                                null; -- label L4833
                                                                -- alt exit (no match)
                                                                b4834 := ("01" = r4822(0 to 1));
                                                                goto_L4836 := b4834;
                                                                if (NOT goto_L4836) then
                                                                  goto_L4842 := (NOT b4834);
                                                                  null; -- label L4842
                                                                  -- alt exit (no match)
                                                                  b4843 := ("10" = r4822(0 to 1));
                                                                  goto_L4845 := b4843;
                                                                  if (NOT goto_L4845) then
                                                                    goto_L4851 := (NOT b4843);
                                                                    null; -- label L4851
                                                                    -- alt exit (no match)
                                                                    -- final pat
                                                                    -- got s@L5 in r4818
                                                                    -- got v'@L4 in r4805
                                                                    r4855 := rewire_setR3_1349(r4818,r4805);
                                                                    statevar0 := r4855;
                                                                    null;
                                                                    goto_L4824 := true;
                                                                  end if;
                                                                  goto_L4824 := goto_L4824;
                                                                  if (NOT goto_L4824) then
                                                                    null; -- label L4845
                                                                    -- got s@L5 in r4818
                                                                    -- got v'@L4 in r4805
                                                                    r4847 := rewire_setR2_1306(r4818,r4805);
                                                                    statevar0 := r4847;
                                                                    null;
                                                                    goto_L4824 := true;
                                                                  end if;
                                                                  goto_L4824 := goto_L4824;
                                                                end if;
                                                                goto_L4824 := goto_L4824;
                                                                if (NOT goto_L4824) then
                                                                  null; -- label L4836
                                                                  -- got s@L5 in r4818
                                                                  -- got v'@L4 in r4805
                                                                  r4838 := rewire_setR1_1262(r4818,r4805);
                                                                  statevar0 := r4838;
                                                                  null;
                                                                  goto_L4824 := true;
                                                                end if;
                                                                goto_L4824 := goto_L4824;
                                                              end if;
                                                              goto_L4824 := goto_L4824;
                                                              if (NOT goto_L4824) then
                                                                null; -- label L4827
                                                                -- got s@L5 in r4818
                                                                -- got v'@L4 in r4805
                                                                r4829 := rewire_setR0_1218(r4818,r4805);
                                                                statevar0 := r4829;
                                                                null;
                                                                goto_L4824 := true;
                                                              end if;
                                                              goto_L4824 := goto_L4824;
                                                              null; -- label L4824
                                                              -- end case
                                                              r4859 := statevar0;
                                                              -- got s@L7 in r4859
                                                              -- got cout@L2 in r4791
                                                              r4863 := rewire_setCFlag_5(r4859,r4791);
                                                              statevar0 := r4863;
                                                              r4866 := statevar0;
                                                              -- got s@L9 in r4866
                                                              -- got v'@L4 in r4805
                                                              r4870 := zeroW8;
                                                              r4872 := eqW8(r4805,r4870);
                                                              r4874 := rewire_setZFlag_48(r4866,r4872);
                                                              statevar0 := r4874;
                                                              r4877 := statevar0;
                                                              -- got s@LB in r4877
                                                              r4880 := rewire_outputs_144(r4877);
                                                              -- got o@LC in r4880
                                                              nextout := r4880;
                                                              state := STATE4885;
                                                              goto_L5439 := true;
                                                            end if;
                                                            goto_L5439 := goto_L5439;
                                                          end if;
                                                          goto_L5439 := goto_L5439;
                                                          if (NOT goto_L5439) then
                                                            null; -- label L4568
                                                            r4567 := statevar0;
                                                            -- got b0@K9 in r4545
                                                            -- got b1@KA in r4547
                                                            r4571 := rewire_mkReg_883(r4545,r4547);
                                                            b4575 := ("00" = r4571(0 to 1));
                                                            goto_L4577 := b4575;
                                                            if (NOT goto_L4577) then
                                                              goto_L4581 := (NOT b4575);
                                                              null; -- label L4581
                                                              -- alt exit (no match)
                                                              b4582 := ("01" = r4571(0 to 1));
                                                              goto_L4584 := b4582;
                                                              if (NOT goto_L4584) then
                                                                goto_L4588 := (NOT b4582);
                                                                null; -- label L4588
                                                                -- alt exit (no match)
                                                                b4589 := ("10" = r4571(0 to 1));
                                                                goto_L4591 := b4589;
                                                                if (NOT goto_L4591) then
                                                                  goto_L4595 := (NOT b4589);
                                                                  null; -- label L4595
                                                                  -- alt exit (no match)
                                                                  -- final pat
                                                                  -- got s@KB in r4567
                                                                  r4598 := rewire_r3_1046(r4567);
                                                                  r4573 := r4598;
                                                                  goto_L4574 := true;
                                                                end if;
                                                                goto_L4574 := goto_L4574;
                                                                if (NOT goto_L4574) then
                                                                  null; -- label L4591
                                                                  -- got s@KB in r4567
                                                                  r4592 := rewire_r2_1008(r4567);
                                                                  r4573 := r4592;
                                                                  goto_L4574 := true;
                                                                end if;
                                                                goto_L4574 := goto_L4574;
                                                              end if;
                                                              goto_L4574 := goto_L4574;
                                                              if (NOT goto_L4574) then
                                                                null; -- label L4584
                                                                -- got s@KB in r4567
                                                                r4585 := rewire_r1_969(r4567);
                                                                r4573 := r4585;
                                                                goto_L4574 := true;
                                                              end if;
                                                              goto_L4574 := goto_L4574;
                                                            end if;
                                                            goto_L4574 := goto_L4574;
                                                            if (NOT goto_L4574) then
                                                              null; -- label L4577
                                                              -- got s@KB in r4567
                                                              r4578 := rewire_r0_930(r4567);
                                                              r4573 := r4578;
                                                              goto_L4574 := true;
                                                            end if;
                                                            goto_L4574 := goto_L4574;
                                                            null; -- label L4574
                                                            -- end case
                                                            -- got v@KC in r4573
                                                            r4602 := oneW8;
                                                            r4604 := "0";
                                                            r4606 := plusCW8(r4573,r4602,r4604);
                                                            -- got p@KD in r4606
                                                            -- final pat
                                                            r4611 := r4606(0 to 0);
                                                            r4613 := r4606(1 to 8);
                                                            b4615 := true;
                                                            b4617 := true;
                                                            -- got x@KE in r4611
                                                            r4609 := r4611;
                                                            -- end case
                                                            -- got p@KD in r4606
                                                            -- final pat
                                                            r4625 := r4606(0 to 0);
                                                            r4627 := r4606(1 to 8);
                                                            b4629 := true;
                                                            b4631 := true;
                                                            -- got x@KG in r4627
                                                            r4623 := r4627;
                                                            -- end case
                                                            r4636 := statevar0;
                                                            -- got b0@K9 in r4545
                                                            -- got b1@KA in r4547
                                                            r4640 := rewire_mkReg_883(r4545,r4547);
                                                            b4643 := ("00" = r4640(0 to 1));
                                                            goto_L4645 := b4643;
                                                            if (NOT goto_L4645) then
                                                              goto_L4651 := (NOT b4643);
                                                              null; -- label L4651
                                                              -- alt exit (no match)
                                                              b4652 := ("01" = r4640(0 to 1));
                                                              goto_L4654 := b4652;
                                                              if (NOT goto_L4654) then
                                                                goto_L4660 := (NOT b4652);
                                                                null; -- label L4660
                                                                -- alt exit (no match)
                                                                b4661 := ("10" = r4640(0 to 1));
                                                                goto_L4663 := b4661;
                                                                if (NOT goto_L4663) then
                                                                  goto_L4669 := (NOT b4661);
                                                                  null; -- label L4669
                                                                  -- alt exit (no match)
                                                                  -- final pat
                                                                  -- got s@KI in r4636
                                                                  -- got v'@KH in r4623
                                                                  r4673 := rewire_setR3_1349(r4636,r4623);
                                                                  statevar0 := r4673;
                                                                  null;
                                                                  goto_L4642 := true;
                                                                end if;
                                                                goto_L4642 := goto_L4642;
                                                                if (NOT goto_L4642) then
                                                                  null; -- label L4663
                                                                  -- got s@KI in r4636
                                                                  -- got v'@KH in r4623
                                                                  r4665 := rewire_setR2_1306(r4636,r4623);
                                                                  statevar0 := r4665;
                                                                  null;
                                                                  goto_L4642 := true;
                                                                end if;
                                                                goto_L4642 := goto_L4642;
                                                              end if;
                                                              goto_L4642 := goto_L4642;
                                                              if (NOT goto_L4642) then
                                                                null; -- label L4654
                                                                -- got s@KI in r4636
                                                                -- got v'@KH in r4623
                                                                r4656 := rewire_setR1_1262(r4636,r4623);
                                                                statevar0 := r4656;
                                                                null;
                                                                goto_L4642 := true;
                                                              end if;
                                                              goto_L4642 := goto_L4642;
                                                            end if;
                                                            goto_L4642 := goto_L4642;
                                                            if (NOT goto_L4642) then
                                                              null; -- label L4645
                                                              -- got s@KI in r4636
                                                              -- got v'@KH in r4623
                                                              r4647 := rewire_setR0_1218(r4636,r4623);
                                                              statevar0 := r4647;
                                                              null;
                                                              goto_L4642 := true;
                                                            end if;
                                                            goto_L4642 := goto_L4642;
                                                            null; -- label L4642
                                                            -- end case
                                                            r4677 := statevar0;
                                                            -- got s@KK in r4677
                                                            -- got cout@KF in r4609
                                                            r4681 := rewire_setCFlag_5(r4677,r4609);
                                                            statevar0 := r4681;
                                                            r4684 := statevar0;
                                                            -- got s@KM in r4684
                                                            -- got v'@KH in r4623
                                                            r4688 := zeroW8;
                                                            r4690 := eqW8(r4623,r4688);
                                                            r4692 := rewire_setZFlag_48(r4684,r4690);
                                                            statevar0 := r4692;
                                                            r4695 := statevar0;
                                                            -- got s@KO in r4695
                                                            r4698 := rewire_outputs_144(r4695);
                                                            -- got o@KP in r4698
                                                            nextout := r4698;
                                                            state := STATE4703;
                                                            goto_L5439 := true;
                                                          end if;
                                                          goto_L5439 := goto_L5439;
                                                        end if;
                                                        goto_L5439 := goto_L5439;
                                                        if (NOT goto_L5439) then
                                                          null; -- label L4469
                                                          r4468 := statevar0;
                                                          -- got b0@K1 in r4446
                                                          -- got b1@K2 in r4448
                                                          r4472 := rewire_mkReg_883(r4446,r4448);
                                                          b4475 := ("00" = r4472(0 to 1));
                                                          goto_L4477 := b4475;
                                                          if (NOT goto_L4477) then
                                                            goto_L4484 := (NOT b4475);
                                                            null; -- label L4484
                                                            -- alt exit (no match)
                                                            b4485 := ("01" = r4472(0 to 1));
                                                            goto_L4487 := b4485;
                                                            if (NOT goto_L4487) then
                                                              goto_L4494 := (NOT b4485);
                                                              null; -- label L4494
                                                              -- alt exit (no match)
                                                              b4495 := ("10" = r4472(0 to 1));
                                                              goto_L4497 := b4495;
                                                              if (NOT goto_L4497) then
                                                                goto_L4504 := (NOT b4495);
                                                                null; -- label L4504
                                                                -- alt exit (no match)
                                                                -- final pat
                                                                -- got s@K3 in r4468
                                                                r4507 := zeroW8;
                                                                r4509 := rewire_setR3_1349(r4468,r4507);
                                                                statevar0 := r4509;
                                                                null;
                                                                goto_L4474 := true;
                                                              end if;
                                                              goto_L4474 := goto_L4474;
                                                              if (NOT goto_L4474) then
                                                                null; -- label L4497
                                                                -- got s@K3 in r4468
                                                                r4498 := zeroW8;
                                                                r4500 := rewire_setR2_1306(r4468,r4498);
                                                                statevar0 := r4500;
                                                                null;
                                                                goto_L4474 := true;
                                                              end if;
                                                              goto_L4474 := goto_L4474;
                                                            end if;
                                                            goto_L4474 := goto_L4474;
                                                            if (NOT goto_L4474) then
                                                              null; -- label L4487
                                                              -- got s@K3 in r4468
                                                              r4488 := zeroW8;
                                                              r4490 := rewire_setR1_1262(r4468,r4488);
                                                              statevar0 := r4490;
                                                              null;
                                                              goto_L4474 := true;
                                                            end if;
                                                            goto_L4474 := goto_L4474;
                                                          end if;
                                                          goto_L4474 := goto_L4474;
                                                          if (NOT goto_L4474) then
                                                            null; -- label L4477
                                                            -- got s@K3 in r4468
                                                            r4478 := zeroW8;
                                                            r4480 := rewire_setR0_1218(r4468,r4478);
                                                            statevar0 := r4480;
                                                            null;
                                                            goto_L4474 := true;
                                                          end if;
                                                          goto_L4474 := goto_L4474;
                                                          null; -- label L4474
                                                          -- end case
                                                          r4513 := statevar0;
                                                          -- got s@K5 in r4513
                                                          r4516 := rewire_outputs_144(r4513);
                                                          -- got o@K6 in r4516
                                                          nextout := r4516;
                                                          state := STATE4521;
                                                          goto_L5439 := true;
                                                        end if;
                                                        goto_L5439 := goto_L5439;
                                                      end if;
                                                      goto_L5439 := goto_L5439;
                                                      if (NOT goto_L5439) then
                                                        null; -- label L4332
                                                        r4331 := statevar0;
                                                        -- got b0@JN in r4309
                                                        -- got b1@JO in r4311
                                                        r4335 := rewire_mkReg_883(r4309,r4311);
                                                        b4339 := ("00" = r4335(0 to 1));
                                                        goto_L4341 := b4339;
                                                        if (NOT goto_L4341) then
                                                          goto_L4345 := (NOT b4339);
                                                          null; -- label L4345
                                                          -- alt exit (no match)
                                                          b4346 := ("01" = r4335(0 to 1));
                                                          goto_L4348 := b4346;
                                                          if (NOT goto_L4348) then
                                                            goto_L4352 := (NOT b4346);
                                                            null; -- label L4352
                                                            -- alt exit (no match)
                                                            b4353 := ("10" = r4335(0 to 1));
                                                            goto_L4355 := b4353;
                                                            if (NOT goto_L4355) then
                                                              goto_L4359 := (NOT b4353);
                                                              null; -- label L4359
                                                              -- alt exit (no match)
                                                              -- final pat
                                                              -- got s@JP in r4331
                                                              r4362 := rewire_r3_1046(r4331);
                                                              r4337 := r4362;
                                                              goto_L4338 := true;
                                                            end if;
                                                            goto_L4338 := goto_L4338;
                                                            if (NOT goto_L4338) then
                                                              null; -- label L4355
                                                              -- got s@JP in r4331
                                                              r4356 := rewire_r2_1008(r4331);
                                                              r4337 := r4356;
                                                              goto_L4338 := true;
                                                            end if;
                                                            goto_L4338 := goto_L4338;
                                                          end if;
                                                          goto_L4338 := goto_L4338;
                                                          if (NOT goto_L4338) then
                                                            null; -- label L4348
                                                            -- got s@JP in r4331
                                                            r4349 := rewire_r1_969(r4331);
                                                            r4337 := r4349;
                                                            goto_L4338 := true;
                                                          end if;
                                                          goto_L4338 := goto_L4338;
                                                        end if;
                                                        goto_L4338 := goto_L4338;
                                                        if (NOT goto_L4338) then
                                                          null; -- label L4341
                                                          -- got s@JP in r4331
                                                          r4342 := rewire_r0_930(r4331);
                                                          r4337 := r4342;
                                                          goto_L4338 := true;
                                                        end if;
                                                        goto_L4338 := goto_L4338;
                                                        null; -- label L4338
                                                        -- end case
                                                        r4365 := statevar0;
                                                        -- got b0@JN in r4309
                                                        -- got b1@JO in r4311
                                                        r4369 := rewire_mkReg_883(r4309,r4311);
                                                        b4372 := ("00" = r4369(0 to 1));
                                                        goto_L4374 := b4372;
                                                        if (NOT goto_L4374) then
                                                          goto_L4382 := (NOT b4372);
                                                          null; -- label L4382
                                                          -- alt exit (no match)
                                                          b4383 := ("01" = r4369(0 to 1));
                                                          goto_L4385 := b4383;
                                                          if (NOT goto_L4385) then
                                                            goto_L4393 := (NOT b4383);
                                                            null; -- label L4393
                                                            -- alt exit (no match)
                                                            b4394 := ("10" = r4369(0 to 1));
                                                            goto_L4396 := b4394;
                                                            if (NOT goto_L4396) then
                                                              goto_L4404 := (NOT b4394);
                                                              null; -- label L4404
                                                              -- alt exit (no match)
                                                              -- final pat
                                                              -- got s@JR in r4365
                                                              -- got v@JQ in r4337
                                                              r4408 := notW8(r4337);
                                                              r4410 := rewire_setR3_1349(r4365,r4408);
                                                              statevar0 := r4410;
                                                              null;
                                                              goto_L4371 := true;
                                                            end if;
                                                            goto_L4371 := goto_L4371;
                                                            if (NOT goto_L4371) then
                                                              null; -- label L4396
                                                              -- got s@JR in r4365
                                                              -- got v@JQ in r4337
                                                              r4398 := notW8(r4337);
                                                              r4400 := rewire_setR2_1306(r4365,r4398);
                                                              statevar0 := r4400;
                                                              null;
                                                              goto_L4371 := true;
                                                            end if;
                                                            goto_L4371 := goto_L4371;
                                                          end if;
                                                          goto_L4371 := goto_L4371;
                                                          if (NOT goto_L4371) then
                                                            null; -- label L4385
                                                            -- got s@JR in r4365
                                                            -- got v@JQ in r4337
                                                            r4387 := notW8(r4337);
                                                            r4389 := rewire_setR1_1262(r4365,r4387);
                                                            statevar0 := r4389;
                                                            null;
                                                            goto_L4371 := true;
                                                          end if;
                                                          goto_L4371 := goto_L4371;
                                                        end if;
                                                        goto_L4371 := goto_L4371;
                                                        if (NOT goto_L4371) then
                                                          null; -- label L4374
                                                          -- got s@JR in r4365
                                                          -- got v@JQ in r4337
                                                          r4376 := notW8(r4337);
                                                          r4378 := rewire_setR0_1218(r4365,r4376);
                                                          statevar0 := r4378;
                                                          null;
                                                          goto_L4371 := true;
                                                        end if;
                                                        goto_L4371 := goto_L4371;
                                                        null; -- label L4371
                                                        -- end case
                                                        r4414 := statevar0;
                                                        -- got s@JT in r4414
                                                        r4417 := rewire_outputs_144(r4414);
                                                        -- got o@JU in r4417
                                                        nextout := r4417;
                                                        state := STATE4422;
                                                        goto_L5439 := true;
                                                      end if;
                                                      goto_L5439 := goto_L5439;
                                                    end if;
                                                    goto_L5439 := goto_L5439;
                                                    if (NOT goto_L5439) then
                                                      null; -- label L4138
                                                      r4137 := statevar0;
                                                      -- got s@J5 in r4137
                                                      r4140 := "1";
                                                      r4142 := rewire_setIEFlag_419(r4137,r4140);
                                                      statevar0 := r4142;
                                                      r4145 := statevar0;
                                                      -- got s@J7 in r4145
                                                      r4180 := rewire_pcSave_4147(r4145);
                                                      r4182 := statevar0;
                                                      -- got s@J9 in r4182
                                                      -- got pc@J8 in r4180
                                                      r4186 := rewire_setPC_1124(r4182,r4180);
                                                      statevar0 := r4186;
                                                      r4189 := statevar0;
                                                      -- got s@JB in r4189
                                                      r4224 := rewire_zsFlag_4191(r4189);
                                                      r4226 := statevar0;
                                                      -- got s@JD in r4226
                                                      -- got z@JC in r4224
                                                      r4230 := rewire_setZFlag_48(r4226,r4224);
                                                      statevar0 := r4230;
                                                      r4233 := statevar0;
                                                      -- got s@JF in r4233
                                                      r4268 := rewire_csFlag_4235(r4233);
                                                      r4270 := statevar0;
                                                      -- got s@JH in r4270
                                                      -- got c@JG in r4268
                                                      r4274 := rewire_setCFlag_5(r4270,r4268);
                                                      statevar0 := r4274;
                                                      r4277 := statevar0;
                                                      -- got s@JJ in r4277
                                                      r4280 := rewire_outputs_144(r4277);
                                                      -- got o@JK in r4280
                                                      nextout := r4280;
                                                      state := STATE4285;
                                                      goto_L5439 := true;
                                                    end if;
                                                    goto_L5439 := goto_L5439;
                                                  end if;
                                                  goto_L5439 := goto_L5439;
                                                  if (NOT goto_L5439) then
                                                    null; -- label L4051
                                                    r4050 := statevar0;
                                                    -- got s@IT in r4050
                                                    r4053 := rewire_outputs_144(r4050);
                                                    r4055 := statevar0;
                                                    -- got s@IV in r4055
                                                    -- got o@IU in r4053
                                                    r4076 := "1";
                                                    r4078 := rewire_setIackOut_4058(r4053,r4076);
                                                    r4080 := rewire_setOutputs_91(r4055,r4078);
                                                    statevar0 := r4080;
                                                    r4083 := statevar0;
                                                    -- got s@J1 in r4083
                                                    r4086 := rewire_outputs_144(r4083);
                                                    -- got o@J2 in r4086
                                                    nextout := r4086;
                                                    state := STATE4091;
                                                    goto_L5439 := true;
                                                  end if;
                                                  goto_L5439 := goto_L5439;
                                                end if;
                                                goto_L5439 := goto_L5439;
                                                if (NOT goto_L5439) then
                                                  null; -- label L3990
                                                  r3989 := statevar0;
                                                  -- got s@IN in r3989
                                                  -- got b0@IM in r3969
                                                  r3993 := rewire_setIEFlag_419(r3989,r3969);
                                                  statevar0 := r3993;
                                                  r3996 := statevar0;
                                                  -- got s@IP in r3996
                                                  r3999 := rewire_outputs_144(r3996);
                                                  -- got o@IQ in r3999
                                                  nextout := r3999;
                                                  state := STATE4004;
                                                  goto_L5439 := true;
                                                end if;
                                                goto_L5439 := goto_L5439;
                                              end if;
                                              goto_L5439 := goto_L5439;
                                              if (NOT goto_L5439) then
                                                null; -- label L3895
                                                r3894 := statevar0;
                                                -- got b0@IC in r3872
                                                -- got b1@ID in r3874
                                                r3898 := rewire_mkReg_883(r3872,r3874);
                                                b3902 := ("00" = r3898(0 to 1));
                                                goto_L3904 := b3902;
                                                if (NOT goto_L3904) then
                                                  goto_L3908 := (NOT b3902);
                                                  null; -- label L3908
                                                  -- alt exit (no match)
                                                  b3909 := ("01" = r3898(0 to 1));
                                                  goto_L3911 := b3909;
                                                  if (NOT goto_L3911) then
                                                    goto_L3915 := (NOT b3909);
                                                    null; -- label L3915
                                                    -- alt exit (no match)
                                                    b3916 := ("10" = r3898(0 to 1));
                                                    goto_L3918 := b3916;
                                                    if (NOT goto_L3918) then
                                                      goto_L3922 := (NOT b3916);
                                                      null; -- label L3922
                                                      -- alt exit (no match)
                                                      -- final pat
                                                      -- got s@IE in r3894
                                                      r3925 := rewire_r3_1046(r3894);
                                                      r3900 := r3925;
                                                      goto_L3901 := true;
                                                    end if;
                                                    goto_L3901 := goto_L3901;
                                                    if (NOT goto_L3901) then
                                                      null; -- label L3918
                                                      -- got s@IE in r3894
                                                      r3919 := rewire_r2_1008(r3894);
                                                      r3900 := r3919;
                                                      goto_L3901 := true;
                                                    end if;
                                                    goto_L3901 := goto_L3901;
                                                  end if;
                                                  goto_L3901 := goto_L3901;
                                                  if (NOT goto_L3901) then
                                                    null; -- label L3911
                                                    -- got s@IE in r3894
                                                    r3912 := rewire_r1_969(r3894);
                                                    r3900 := r3912;
                                                    goto_L3901 := true;
                                                  end if;
                                                  goto_L3901 := goto_L3901;
                                                end if;
                                                goto_L3901 := goto_L3901;
                                                if (NOT goto_L3901) then
                                                  null; -- label L3904
                                                  -- got s@IE in r3894
                                                  r3905 := rewire_r0_930(r3894);
                                                  r3900 := r3905;
                                                  goto_L3901 := true;
                                                end if;
                                                goto_L3901 := goto_L3901;
                                                null; -- label L3901
                                                -- end case
                                                r3928 := statevar0;
                                                -- got s@IG in r3928
                                                -- got a@IF in r3900
                                                r3932 := rewire_setPC_1124(r3928,r3900);
                                                statevar0 := r3932;
                                                r3935 := statevar0;
                                                -- got s@II in r3935
                                                r3938 := rewire_outputs_144(r3935);
                                                -- got o@IJ in r3938
                                                nextout := r3938;
                                                state := STATE3943;
                                                goto_L5439 := true;
                                              end if;
                                              goto_L5439 := goto_L5439;
                                            end if;
                                            goto_L5439 := goto_L5439;
                                            if (NOT goto_L5439) then
                                              null; -- label L3784
                                              r3783 := statevar0;
                                              -- got s@I2 in r3783
                                              r3786 := rewire_cFlag_536(r3783);
                                              -- got c@I3 in r3786
                                              r3789 := notBit(r3786);
                                              b3792 := ("1" = r3789(0 to 0));
                                              goto_L3795 := b3792;
                                              if (NOT goto_L3795) then
                                                goto_L3836 := (NOT b3792);
                                                null; -- label L3836
                                                -- alt exit (no match)
                                                -- final pat
                                                null;
                                                null;
                                                goto_L3791 := true;
                                              end if;
                                              goto_L3791 := goto_L3791;
                                              if (NOT goto_L3791) then
                                                null; -- label L3795
                                                r3794 := statevar0;
                                                -- got b0@I0 in r3761
                                                -- got b1@I1 in r3763
                                                r3798 := rewire_mkReg_883(r3761,r3763);
                                                b3802 := ("00" = r3798(0 to 1));
                                                goto_L3804 := b3802;
                                                if (NOT goto_L3804) then
                                                  goto_L3808 := (NOT b3802);
                                                  null; -- label L3808
                                                  -- alt exit (no match)
                                                  b3809 := ("01" = r3798(0 to 1));
                                                  goto_L3811 := b3809;
                                                  if (NOT goto_L3811) then
                                                    goto_L3815 := (NOT b3809);
                                                    null; -- label L3815
                                                    -- alt exit (no match)
                                                    b3816 := ("10" = r3798(0 to 1));
                                                    goto_L3818 := b3816;
                                                    if (NOT goto_L3818) then
                                                      goto_L3822 := (NOT b3816);
                                                      null; -- label L3822
                                                      -- alt exit (no match)
                                                      -- final pat
                                                      -- got s@I4 in r3794
                                                      r3825 := rewire_r3_1046(r3794);
                                                      r3800 := r3825;
                                                      goto_L3801 := true;
                                                    end if;
                                                    goto_L3801 := goto_L3801;
                                                    if (NOT goto_L3801) then
                                                      null; -- label L3818
                                                      -- got s@I4 in r3794
                                                      r3819 := rewire_r2_1008(r3794);
                                                      r3800 := r3819;
                                                      goto_L3801 := true;
                                                    end if;
                                                    goto_L3801 := goto_L3801;
                                                  end if;
                                                  goto_L3801 := goto_L3801;
                                                  if (NOT goto_L3801) then
                                                    null; -- label L3811
                                                    -- got s@I4 in r3794
                                                    r3812 := rewire_r1_969(r3794);
                                                    r3800 := r3812;
                                                    goto_L3801 := true;
                                                  end if;
                                                  goto_L3801 := goto_L3801;
                                                end if;
                                                goto_L3801 := goto_L3801;
                                                if (NOT goto_L3801) then
                                                  null; -- label L3804
                                                  -- got s@I4 in r3794
                                                  r3805 := rewire_r0_930(r3794);
                                                  r3800 := r3805;
                                                  goto_L3801 := true;
                                                end if;
                                                goto_L3801 := goto_L3801;
                                                null; -- label L3801
                                                -- end case
                                                r3828 := statevar0;
                                                -- got s@I6 in r3828
                                                -- got a@I5 in r3800
                                                r3832 := rewire_setPC_1124(r3828,r3800);
                                                statevar0 := r3832;
                                                null;
                                                goto_L3791 := true;
                                              end if;
                                              goto_L3791 := goto_L3791;
                                              null; -- label L3791
                                              -- end case
                                              r3840 := statevar0;
                                              -- got s@I8 in r3840
                                              r3843 := rewire_outputs_144(r3840);
                                              -- got o@I9 in r3843
                                              nextout := r3843;
                                              state := STATE3848;
                                              goto_L5439 := true;
                                            end if;
                                            goto_L5439 := goto_L5439;
                                          end if;
                                          goto_L5439 := goto_L5439;
                                          if (NOT goto_L5439) then
                                            null; -- label L3675
                                            r3674 := statevar0;
                                            -- got s@HM in r3674
                                            r3677 := rewire_cFlag_536(r3674);
                                            -- got c@HN in r3677
                                            b3681 := ("1" = r3677(0 to 0));
                                            goto_L3684 := b3681;
                                            if (NOT goto_L3684) then
                                              goto_L3725 := (NOT b3681);
                                              null; -- label L3725
                                              -- alt exit (no match)
                                              -- final pat
                                              null;
                                              null;
                                              goto_L3680 := true;
                                            end if;
                                            goto_L3680 := goto_L3680;
                                            if (NOT goto_L3680) then
                                              null; -- label L3684
                                              r3683 := statevar0;
                                              -- got b0@HK in r3652
                                              -- got b1@HL in r3654
                                              r3687 := rewire_mkReg_883(r3652,r3654);
                                              b3691 := ("00" = r3687(0 to 1));
                                              goto_L3693 := b3691;
                                              if (NOT goto_L3693) then
                                                goto_L3697 := (NOT b3691);
                                                null; -- label L3697
                                                -- alt exit (no match)
                                                b3698 := ("01" = r3687(0 to 1));
                                                goto_L3700 := b3698;
                                                if (NOT goto_L3700) then
                                                  goto_L3704 := (NOT b3698);
                                                  null; -- label L3704
                                                  -- alt exit (no match)
                                                  b3705 := ("10" = r3687(0 to 1));
                                                  goto_L3707 := b3705;
                                                  if (NOT goto_L3707) then
                                                    goto_L3711 := (NOT b3705);
                                                    null; -- label L3711
                                                    -- alt exit (no match)
                                                    -- final pat
                                                    -- got s@HO in r3683
                                                    r3714 := rewire_r3_1046(r3683);
                                                    r3689 := r3714;
                                                    goto_L3690 := true;
                                                  end if;
                                                  goto_L3690 := goto_L3690;
                                                  if (NOT goto_L3690) then
                                                    null; -- label L3707
                                                    -- got s@HO in r3683
                                                    r3708 := rewire_r2_1008(r3683);
                                                    r3689 := r3708;
                                                    goto_L3690 := true;
                                                  end if;
                                                  goto_L3690 := goto_L3690;
                                                end if;
                                                goto_L3690 := goto_L3690;
                                                if (NOT goto_L3690) then
                                                  null; -- label L3700
                                                  -- got s@HO in r3683
                                                  r3701 := rewire_r1_969(r3683);
                                                  r3689 := r3701;
                                                  goto_L3690 := true;
                                                end if;
                                                goto_L3690 := goto_L3690;
                                              end if;
                                              goto_L3690 := goto_L3690;
                                              if (NOT goto_L3690) then
                                                null; -- label L3693
                                                -- got s@HO in r3683
                                                r3694 := rewire_r0_930(r3683);
                                                r3689 := r3694;
                                                goto_L3690 := true;
                                              end if;
                                              goto_L3690 := goto_L3690;
                                              null; -- label L3690
                                              -- end case
                                              r3717 := statevar0;
                                              -- got s@HQ in r3717
                                              -- got a@HP in r3689
                                              r3721 := rewire_setPC_1124(r3717,r3689);
                                              statevar0 := r3721;
                                              null;
                                              goto_L3680 := true;
                                            end if;
                                            goto_L3680 := goto_L3680;
                                            null; -- label L3680
                                            -- end case
                                            r3729 := statevar0;
                                            -- got s@HS in r3729
                                            r3732 := rewire_outputs_144(r3729);
                                            -- got o@HT in r3732
                                            nextout := r3732;
                                            state := STATE3737;
                                            goto_L5439 := true;
                                          end if;
                                          goto_L5439 := goto_L5439;
                                        end if;
                                        goto_L5439 := goto_L5439;
                                        if (NOT goto_L5439) then
                                          null; -- label L3564
                                          r3563 := statevar0;
                                          -- got s@HA in r3563
                                          r3566 := rewire_zFlag_499(r3563);
                                          -- got z@HB in r3566
                                          r3569 := notBit(r3566);
                                          b3572 := ("1" = r3569(0 to 0));
                                          goto_L3575 := b3572;
                                          if (NOT goto_L3575) then
                                            goto_L3616 := (NOT b3572);
                                            null; -- label L3616
                                            -- alt exit (no match)
                                            -- final pat
                                            null;
                                            null;
                                            goto_L3571 := true;
                                          end if;
                                          goto_L3571 := goto_L3571;
                                          if (NOT goto_L3571) then
                                            null; -- label L3575
                                            r3574 := statevar0;
                                            -- got b0@H8 in r3541
                                            -- got b1@H9 in r3543
                                            r3578 := rewire_mkReg_883(r3541,r3543);
                                            b3582 := ("00" = r3578(0 to 1));
                                            goto_L3584 := b3582;
                                            if (NOT goto_L3584) then
                                              goto_L3588 := (NOT b3582);
                                              null; -- label L3588
                                              -- alt exit (no match)
                                              b3589 := ("01" = r3578(0 to 1));
                                              goto_L3591 := b3589;
                                              if (NOT goto_L3591) then
                                                goto_L3595 := (NOT b3589);
                                                null; -- label L3595
                                                -- alt exit (no match)
                                                b3596 := ("10" = r3578(0 to 1));
                                                goto_L3598 := b3596;
                                                if (NOT goto_L3598) then
                                                  goto_L3602 := (NOT b3596);
                                                  null; -- label L3602
                                                  -- alt exit (no match)
                                                  -- final pat
                                                  -- got s@HC in r3574
                                                  r3605 := rewire_r3_1046(r3574);
                                                  r3580 := r3605;
                                                  goto_L3581 := true;
                                                end if;
                                                goto_L3581 := goto_L3581;
                                                if (NOT goto_L3581) then
                                                  null; -- label L3598
                                                  -- got s@HC in r3574
                                                  r3599 := rewire_r2_1008(r3574);
                                                  r3580 := r3599;
                                                  goto_L3581 := true;
                                                end if;
                                                goto_L3581 := goto_L3581;
                                              end if;
                                              goto_L3581 := goto_L3581;
                                              if (NOT goto_L3581) then
                                                null; -- label L3591
                                                -- got s@HC in r3574
                                                r3592 := rewire_r1_969(r3574);
                                                r3580 := r3592;
                                                goto_L3581 := true;
                                              end if;
                                              goto_L3581 := goto_L3581;
                                            end if;
                                            goto_L3581 := goto_L3581;
                                            if (NOT goto_L3581) then
                                              null; -- label L3584
                                              -- got s@HC in r3574
                                              r3585 := rewire_r0_930(r3574);
                                              r3580 := r3585;
                                              goto_L3581 := true;
                                            end if;
                                            goto_L3581 := goto_L3581;
                                            null; -- label L3581
                                            -- end case
                                            r3608 := statevar0;
                                            -- got s@HE in r3608
                                            -- got a@HD in r3580
                                            r3612 := rewire_setPC_1124(r3608,r3580);
                                            statevar0 := r3612;
                                            null;
                                            goto_L3571 := true;
                                          end if;
                                          goto_L3571 := goto_L3571;
                                          null; -- label L3571
                                          -- end case
                                          r3620 := statevar0;
                                          -- got s@HG in r3620
                                          r3623 := rewire_outputs_144(r3620);
                                          -- got o@HH in r3623
                                          nextout := r3623;
                                          state := STATE3628;
                                          goto_L5439 := true;
                                        end if;
                                        goto_L5439 := goto_L5439;
                                      end if;
                                      goto_L5439 := goto_L5439;
                                      if (NOT goto_L5439) then
                                        null; -- label L3455
                                        r3454 := statevar0;
                                        -- got s@GU in r3454
                                        r3457 := rewire_zFlag_499(r3454);
                                        -- got z@GV in r3457
                                        b3461 := ("1" = r3457(0 to 0));
                                        goto_L3464 := b3461;
                                        if (NOT goto_L3464) then
                                          goto_L3505 := (NOT b3461);
                                          null; -- label L3505
                                          -- alt exit (no match)
                                          -- final pat
                                          null;
                                          null;
                                          goto_L3460 := true;
                                        end if;
                                        goto_L3460 := goto_L3460;
                                        if (NOT goto_L3460) then
                                          null; -- label L3464
                                          r3463 := statevar0;
                                          -- got b0@GS in r3432
                                          -- got b1@GT in r3434
                                          r3467 := rewire_mkReg_883(r3432,r3434);
                                          b3471 := ("00" = r3467(0 to 1));
                                          goto_L3473 := b3471;
                                          if (NOT goto_L3473) then
                                            goto_L3477 := (NOT b3471);
                                            null; -- label L3477
                                            -- alt exit (no match)
                                            b3478 := ("01" = r3467(0 to 1));
                                            goto_L3480 := b3478;
                                            if (NOT goto_L3480) then
                                              goto_L3484 := (NOT b3478);
                                              null; -- label L3484
                                              -- alt exit (no match)
                                              b3485 := ("10" = r3467(0 to 1));
                                              goto_L3487 := b3485;
                                              if (NOT goto_L3487) then
                                                goto_L3491 := (NOT b3485);
                                                null; -- label L3491
                                                -- alt exit (no match)
                                                -- final pat
                                                -- got s@H0 in r3463
                                                r3494 := rewire_r3_1046(r3463);
                                                r3469 := r3494;
                                                goto_L3470 := true;
                                              end if;
                                              goto_L3470 := goto_L3470;
                                              if (NOT goto_L3470) then
                                                null; -- label L3487
                                                -- got s@H0 in r3463
                                                r3488 := rewire_r2_1008(r3463);
                                                r3469 := r3488;
                                                goto_L3470 := true;
                                              end if;
                                              goto_L3470 := goto_L3470;
                                            end if;
                                            goto_L3470 := goto_L3470;
                                            if (NOT goto_L3470) then
                                              null; -- label L3480
                                              -- got s@H0 in r3463
                                              r3481 := rewire_r1_969(r3463);
                                              r3469 := r3481;
                                              goto_L3470 := true;
                                            end if;
                                            goto_L3470 := goto_L3470;
                                          end if;
                                          goto_L3470 := goto_L3470;
                                          if (NOT goto_L3470) then
                                            null; -- label L3473
                                            -- got s@H0 in r3463
                                            r3474 := rewire_r0_930(r3463);
                                            r3469 := r3474;
                                            goto_L3470 := true;
                                          end if;
                                          goto_L3470 := goto_L3470;
                                          null; -- label L3470
                                          -- end case
                                          r3497 := statevar0;
                                          -- got s@H2 in r3497
                                          -- got a@H1 in r3469
                                          r3501 := rewire_setPC_1124(r3497,r3469);
                                          statevar0 := r3501;
                                          null;
                                          goto_L3460 := true;
                                        end if;
                                        goto_L3460 := goto_L3460;
                                        null; -- label L3460
                                        -- end case
                                        r3509 := statevar0;
                                        -- got s@H4 in r3509
                                        r3512 := rewire_outputs_144(r3509);
                                        -- got o@H5 in r3512
                                        nextout := r3512;
                                        state := STATE3517;
                                        goto_L5439 := true;
                                      end if;
                                      goto_L5439 := goto_L5439;
                                    end if;
                                    goto_L5439 := goto_L5439;
                                    if (NOT goto_L5439) then
                                      null; -- label L3281
                                      r3280 := statevar0;
                                      -- got b0@G7 in r3254
                                      -- got b1@G8 in r3256
                                      r3284 := rewire_mkReg_883(r3254,r3256);
                                      b3288 := ("00" = r3284(0 to 1));
                                      goto_L3290 := b3288;
                                      if (NOT goto_L3290) then
                                        goto_L3294 := (NOT b3288);
                                        null; -- label L3294
                                        -- alt exit (no match)
                                        b3295 := ("01" = r3284(0 to 1));
                                        goto_L3297 := b3295;
                                        if (NOT goto_L3297) then
                                          goto_L3301 := (NOT b3295);
                                          null; -- label L3301
                                          -- alt exit (no match)
                                          b3302 := ("10" = r3284(0 to 1));
                                          goto_L3304 := b3302;
                                          if (NOT goto_L3304) then
                                            goto_L3308 := (NOT b3302);
                                            null; -- label L3308
                                            -- alt exit (no match)
                                            -- final pat
                                            -- got s@GB in r3280
                                            r3311 := rewire_r3_1046(r3280);
                                            r3286 := r3311;
                                            goto_L3287 := true;
                                          end if;
                                          goto_L3287 := goto_L3287;
                                          if (NOT goto_L3287) then
                                            null; -- label L3304
                                            -- got s@GB in r3280
                                            r3305 := rewire_r2_1008(r3280);
                                            r3286 := r3305;
                                            goto_L3287 := true;
                                          end if;
                                          goto_L3287 := goto_L3287;
                                        end if;
                                        goto_L3287 := goto_L3287;
                                        if (NOT goto_L3287) then
                                          null; -- label L3297
                                          -- got s@GB in r3280
                                          r3298 := rewire_r1_969(r3280);
                                          r3286 := r3298;
                                          goto_L3287 := true;
                                        end if;
                                        goto_L3287 := goto_L3287;
                                      end if;
                                      goto_L3287 := goto_L3287;
                                      if (NOT goto_L3287) then
                                        null; -- label L3290
                                        -- got s@GB in r3280
                                        r3291 := rewire_r0_930(r3280);
                                        r3286 := r3291;
                                        goto_L3287 := true;
                                      end if;
                                      goto_L3287 := goto_L3287;
                                      null; -- label L3287
                                      -- end case
                                      r3314 := statevar0;
                                      -- got c0@G9 in r3258
                                      -- got c1@GA in r3260
                                      r3318 := rewire_mkReg_883(r3258,r3260);
                                      b3322 := ("00" = r3318(0 to 1));
                                      goto_L3324 := b3322;
                                      if (NOT goto_L3324) then
                                        goto_L3328 := (NOT b3322);
                                        null; -- label L3328
                                        -- alt exit (no match)
                                        b3329 := ("01" = r3318(0 to 1));
                                        goto_L3331 := b3329;
                                        if (NOT goto_L3331) then
                                          goto_L3335 := (NOT b3329);
                                          null; -- label L3335
                                          -- alt exit (no match)
                                          b3336 := ("10" = r3318(0 to 1));
                                          goto_L3338 := b3336;
                                          if (NOT goto_L3338) then
                                            goto_L3342 := (NOT b3336);
                                            null; -- label L3342
                                            -- alt exit (no match)
                                            -- final pat
                                            -- got s@GD in r3314
                                            r3345 := rewire_r3_1046(r3314);
                                            r3320 := r3345;
                                            goto_L3321 := true;
                                          end if;
                                          goto_L3321 := goto_L3321;
                                          if (NOT goto_L3321) then
                                            null; -- label L3338
                                            -- got s@GD in r3314
                                            r3339 := rewire_r2_1008(r3314);
                                            r3320 := r3339;
                                            goto_L3321 := true;
                                          end if;
                                          goto_L3321 := goto_L3321;
                                        end if;
                                        goto_L3321 := goto_L3321;
                                        if (NOT goto_L3321) then
                                          null; -- label L3331
                                          -- got s@GD in r3314
                                          r3332 := rewire_r1_969(r3314);
                                          r3320 := r3332;
                                          goto_L3321 := true;
                                        end if;
                                        goto_L3321 := goto_L3321;
                                      end if;
                                      goto_L3321 := goto_L3321;
                                      if (NOT goto_L3321) then
                                        null; -- label L3324
                                        -- got s@GD in r3314
                                        r3325 := rewire_r0_930(r3314);
                                        r3320 := r3325;
                                        goto_L3321 := true;
                                      end if;
                                      goto_L3321 := goto_L3321;
                                      null; -- label L3321
                                      -- end case
                                      -- got vD@GC in r3286
                                      -- got vS@GE in r3320
                                      r3350 := "0";
                                      r3352 := minusCW8(r3286,r3320,r3350);
                                      -- got p@GF in r3352
                                      -- final pat
                                      r3357 := r3352(0 to 0);
                                      r3359 := r3352(1 to 8);
                                      b3361 := true;
                                      b3363 := true;
                                      -- got x@GG in r3357
                                      r3355 := r3357;
                                      -- end case
                                      -- got p@GF in r3352
                                      -- final pat
                                      r3371 := r3352(0 to 0);
                                      r3373 := r3352(1 to 8);
                                      b3375 := true;
                                      b3377 := true;
                                      -- got x@GI in r3373
                                      r3369 := r3373;
                                      -- end case
                                      r3382 := statevar0;
                                      -- got s@GK in r3382
                                      -- got c@GH in r3355
                                      r3386 := rewire_setCFlag_5(r3382,r3355);
                                      statevar0 := r3386;
                                      r3389 := statevar0;
                                      -- got s@GM in r3389
                                      -- got r@GJ in r3369
                                      r3393 := zeroW8;
                                      r3395 := eqW8(r3369,r3393);
                                      r3397 := rewire_setZFlag_48(r3389,r3395);
                                      statevar0 := r3397;
                                      r3400 := statevar0;
                                      -- got s@GO in r3400
                                      r3403 := rewire_outputs_144(r3400);
                                      -- got o@GP in r3403
                                      nextout := r3403;
                                      state := STATE3408;
                                      goto_L5439 := true;
                                    end if;
                                    goto_L5439 := goto_L5439;
                                  end if;
                                  goto_L5439 := goto_L5439;
                                  if (NOT goto_L5439) then
                                    null; -- label L3095
                                    r3094 := statevar0;
                                    -- got b0@FK in r3068
                                    -- got b1@FL in r3070
                                    r3098 := rewire_mkReg_883(r3068,r3070);
                                    b3102 := ("00" = r3098(0 to 1));
                                    goto_L3104 := b3102;
                                    if (NOT goto_L3104) then
                                      goto_L3108 := (NOT b3102);
                                      null; -- label L3108
                                      -- alt exit (no match)
                                      b3109 := ("01" = r3098(0 to 1));
                                      goto_L3111 := b3109;
                                      if (NOT goto_L3111) then
                                        goto_L3115 := (NOT b3109);
                                        null; -- label L3115
                                        -- alt exit (no match)
                                        b3116 := ("10" = r3098(0 to 1));
                                        goto_L3118 := b3116;
                                        if (NOT goto_L3118) then
                                          goto_L3122 := (NOT b3116);
                                          null; -- label L3122
                                          -- alt exit (no match)
                                          -- final pat
                                          -- got s@FO in r3094
                                          r3125 := rewire_r3_1046(r3094);
                                          r3100 := r3125;
                                          goto_L3101 := true;
                                        end if;
                                        goto_L3101 := goto_L3101;
                                        if (NOT goto_L3101) then
                                          null; -- label L3118
                                          -- got s@FO in r3094
                                          r3119 := rewire_r2_1008(r3094);
                                          r3100 := r3119;
                                          goto_L3101 := true;
                                        end if;
                                        goto_L3101 := goto_L3101;
                                      end if;
                                      goto_L3101 := goto_L3101;
                                      if (NOT goto_L3101) then
                                        null; -- label L3111
                                        -- got s@FO in r3094
                                        r3112 := rewire_r1_969(r3094);
                                        r3100 := r3112;
                                        goto_L3101 := true;
                                      end if;
                                      goto_L3101 := goto_L3101;
                                    end if;
                                    goto_L3101 := goto_L3101;
                                    if (NOT goto_L3101) then
                                      null; -- label L3104
                                      -- got s@FO in r3094
                                      r3105 := rewire_r0_930(r3094);
                                      r3100 := r3105;
                                      goto_L3101 := true;
                                    end if;
                                    goto_L3101 := goto_L3101;
                                    null; -- label L3101
                                    -- end case
                                    r3128 := statevar0;
                                    -- got c0@FM in r3072
                                    -- got c1@FN in r3074
                                    r3132 := rewire_mkReg_883(r3072,r3074);
                                    b3136 := ("00" = r3132(0 to 1));
                                    goto_L3138 := b3136;
                                    if (NOT goto_L3138) then
                                      goto_L3142 := (NOT b3136);
                                      null; -- label L3142
                                      -- alt exit (no match)
                                      b3143 := ("01" = r3132(0 to 1));
                                      goto_L3145 := b3143;
                                      if (NOT goto_L3145) then
                                        goto_L3149 := (NOT b3143);
                                        null; -- label L3149
                                        -- alt exit (no match)
                                        b3150 := ("10" = r3132(0 to 1));
                                        goto_L3152 := b3150;
                                        if (NOT goto_L3152) then
                                          goto_L3156 := (NOT b3150);
                                          null; -- label L3156
                                          -- alt exit (no match)
                                          -- final pat
                                          -- got s@FQ in r3128
                                          r3159 := rewire_r3_1046(r3128);
                                          r3134 := r3159;
                                          goto_L3135 := true;
                                        end if;
                                        goto_L3135 := goto_L3135;
                                        if (NOT goto_L3135) then
                                          null; -- label L3152
                                          -- got s@FQ in r3128
                                          r3153 := rewire_r2_1008(r3128);
                                          r3134 := r3153;
                                          goto_L3135 := true;
                                        end if;
                                        goto_L3135 := goto_L3135;
                                      end if;
                                      goto_L3135 := goto_L3135;
                                      if (NOT goto_L3135) then
                                        null; -- label L3145
                                        -- got s@FQ in r3128
                                        r3146 := rewire_r1_969(r3128);
                                        r3134 := r3146;
                                        goto_L3135 := true;
                                      end if;
                                      goto_L3135 := goto_L3135;
                                    end if;
                                    goto_L3135 := goto_L3135;
                                    if (NOT goto_L3135) then
                                      null; -- label L3138
                                      -- got s@FQ in r3128
                                      r3139 := rewire_r0_930(r3128);
                                      r3134 := r3139;
                                      goto_L3135 := true;
                                    end if;
                                    goto_L3135 := goto_L3135;
                                    null; -- label L3135
                                    -- end case
                                    -- got vD@FP in r3100
                                    -- got vS@FR in r3134
                                    r3164 := xorW8(r3100,r3134);
                                    r3166 := statevar0;
                                    -- got b0@FK in r3068
                                    -- got b1@FL in r3070
                                    r3170 := rewire_mkReg_883(r3068,r3070);
                                    b3173 := ("00" = r3170(0 to 1));
                                    goto_L3175 := b3173;
                                    if (NOT goto_L3175) then
                                      goto_L3181 := (NOT b3173);
                                      null; -- label L3181
                                      -- alt exit (no match)
                                      b3182 := ("01" = r3170(0 to 1));
                                      goto_L3184 := b3182;
                                      if (NOT goto_L3184) then
                                        goto_L3190 := (NOT b3182);
                                        null; -- label L3190
                                        -- alt exit (no match)
                                        b3191 := ("10" = r3170(0 to 1));
                                        goto_L3193 := b3191;
                                        if (NOT goto_L3193) then
                                          goto_L3199 := (NOT b3191);
                                          null; -- label L3199
                                          -- alt exit (no match)
                                          -- final pat
                                          -- got s@FT in r3166
                                          -- got vD'@FS in r3164
                                          r3203 := rewire_setR3_1349(r3166,r3164);
                                          statevar0 := r3203;
                                          null;
                                          goto_L3172 := true;
                                        end if;
                                        goto_L3172 := goto_L3172;
                                        if (NOT goto_L3172) then
                                          null; -- label L3193
                                          -- got s@FT in r3166
                                          -- got vD'@FS in r3164
                                          r3195 := rewire_setR2_1306(r3166,r3164);
                                          statevar0 := r3195;
                                          null;
                                          goto_L3172 := true;
                                        end if;
                                        goto_L3172 := goto_L3172;
                                      end if;
                                      goto_L3172 := goto_L3172;
                                      if (NOT goto_L3172) then
                                        null; -- label L3184
                                        -- got s@FT in r3166
                                        -- got vD'@FS in r3164
                                        r3186 := rewire_setR1_1262(r3166,r3164);
                                        statevar0 := r3186;
                                        null;
                                        goto_L3172 := true;
                                      end if;
                                      goto_L3172 := goto_L3172;
                                    end if;
                                    goto_L3172 := goto_L3172;
                                    if (NOT goto_L3172) then
                                      null; -- label L3175
                                      -- got s@FT in r3166
                                      -- got vD'@FS in r3164
                                      r3177 := rewire_setR0_1218(r3166,r3164);
                                      statevar0 := r3177;
                                      null;
                                      goto_L3172 := true;
                                    end if;
                                    goto_L3172 := goto_L3172;
                                    null; -- label L3172
                                    -- end case
                                    r3207 := statevar0;
                                    -- got s@FV in r3207
                                    r3210 := "0";
                                    r3212 := rewire_setCFlag_5(r3207,r3210);
                                    statevar0 := r3212;
                                    r3215 := statevar0;
                                    -- got s@G1 in r3215
                                    -- got vD'@FS in r3164
                                    r3219 := zeroW8;
                                    r3221 := eqW8(r3164,r3219);
                                    r3223 := rewire_setZFlag_48(r3215,r3221);
                                    statevar0 := r3223;
                                    r3226 := statevar0;
                                    -- got s@G3 in r3226
                                    r3229 := rewire_outputs_144(r3226);
                                    -- got o@G4 in r3229
                                    nextout := r3229;
                                    state := STATE3234;
                                    goto_L5439 := true;
                                  end if;
                                  goto_L5439 := goto_L5439;
                                end if;
                                goto_L5439 := goto_L5439;
                                if (NOT goto_L5439) then
                                  null; -- label L2909
                                  r2908 := statevar0;
                                  -- got b0@F1 in r2882
                                  -- got b1@F2 in r2884
                                  r2912 := rewire_mkReg_883(r2882,r2884);
                                  b2916 := ("00" = r2912(0 to 1));
                                  goto_L2918 := b2916;
                                  if (NOT goto_L2918) then
                                    goto_L2922 := (NOT b2916);
                                    null; -- label L2922
                                    -- alt exit (no match)
                                    b2923 := ("01" = r2912(0 to 1));
                                    goto_L2925 := b2923;
                                    if (NOT goto_L2925) then
                                      goto_L2929 := (NOT b2923);
                                      null; -- label L2929
                                      -- alt exit (no match)
                                      b2930 := ("10" = r2912(0 to 1));
                                      goto_L2932 := b2930;
                                      if (NOT goto_L2932) then
                                        goto_L2936 := (NOT b2930);
                                        null; -- label L2936
                                        -- alt exit (no match)
                                        -- final pat
                                        -- got s@F5 in r2908
                                        r2939 := rewire_r3_1046(r2908);
                                        r2914 := r2939;
                                        goto_L2915 := true;
                                      end if;
                                      goto_L2915 := goto_L2915;
                                      if (NOT goto_L2915) then
                                        null; -- label L2932
                                        -- got s@F5 in r2908
                                        r2933 := rewire_r2_1008(r2908);
                                        r2914 := r2933;
                                        goto_L2915 := true;
                                      end if;
                                      goto_L2915 := goto_L2915;
                                    end if;
                                    goto_L2915 := goto_L2915;
                                    if (NOT goto_L2915) then
                                      null; -- label L2925
                                      -- got s@F5 in r2908
                                      r2926 := rewire_r1_969(r2908);
                                      r2914 := r2926;
                                      goto_L2915 := true;
                                    end if;
                                    goto_L2915 := goto_L2915;
                                  end if;
                                  goto_L2915 := goto_L2915;
                                  if (NOT goto_L2915) then
                                    null; -- label L2918
                                    -- got s@F5 in r2908
                                    r2919 := rewire_r0_930(r2908);
                                    r2914 := r2919;
                                    goto_L2915 := true;
                                  end if;
                                  goto_L2915 := goto_L2915;
                                  null; -- label L2915
                                  -- end case
                                  r2942 := statevar0;
                                  -- got c0@F3 in r2886
                                  -- got c1@F4 in r2888
                                  r2946 := rewire_mkReg_883(r2886,r2888);
                                  b2950 := ("00" = r2946(0 to 1));
                                  goto_L2952 := b2950;
                                  if (NOT goto_L2952) then
                                    goto_L2956 := (NOT b2950);
                                    null; -- label L2956
                                    -- alt exit (no match)
                                    b2957 := ("01" = r2946(0 to 1));
                                    goto_L2959 := b2957;
                                    if (NOT goto_L2959) then
                                      goto_L2963 := (NOT b2957);
                                      null; -- label L2963
                                      -- alt exit (no match)
                                      b2964 := ("10" = r2946(0 to 1));
                                      goto_L2966 := b2964;
                                      if (NOT goto_L2966) then
                                        goto_L2970 := (NOT b2964);
                                        null; -- label L2970
                                        -- alt exit (no match)
                                        -- final pat
                                        -- got s@F7 in r2942
                                        r2973 := rewire_r3_1046(r2942);
                                        r2948 := r2973;
                                        goto_L2949 := true;
                                      end if;
                                      goto_L2949 := goto_L2949;
                                      if (NOT goto_L2949) then
                                        null; -- label L2966
                                        -- got s@F7 in r2942
                                        r2967 := rewire_r2_1008(r2942);
                                        r2948 := r2967;
                                        goto_L2949 := true;
                                      end if;
                                      goto_L2949 := goto_L2949;
                                    end if;
                                    goto_L2949 := goto_L2949;
                                    if (NOT goto_L2949) then
                                      null; -- label L2959
                                      -- got s@F7 in r2942
                                      r2960 := rewire_r1_969(r2942);
                                      r2948 := r2960;
                                      goto_L2949 := true;
                                    end if;
                                    goto_L2949 := goto_L2949;
                                  end if;
                                  goto_L2949 := goto_L2949;
                                  if (NOT goto_L2949) then
                                    null; -- label L2952
                                    -- got s@F7 in r2942
                                    r2953 := rewire_r0_930(r2942);
                                    r2948 := r2953;
                                    goto_L2949 := true;
                                  end if;
                                  goto_L2949 := goto_L2949;
                                  null; -- label L2949
                                  -- end case
                                  -- got vD@F6 in r2914
                                  -- got vS@F8 in r2948
                                  r2978 := andW8(r2914,r2948);
                                  r2980 := statevar0;
                                  -- got b0@F1 in r2882
                                  -- got b1@F2 in r2884
                                  r2984 := rewire_mkReg_883(r2882,r2884);
                                  b2987 := ("00" = r2984(0 to 1));
                                  goto_L2989 := b2987;
                                  if (NOT goto_L2989) then
                                    goto_L2995 := (NOT b2987);
                                    null; -- label L2995
                                    -- alt exit (no match)
                                    b2996 := ("01" = r2984(0 to 1));
                                    goto_L2998 := b2996;
                                    if (NOT goto_L2998) then
                                      goto_L3004 := (NOT b2996);
                                      null; -- label L3004
                                      -- alt exit (no match)
                                      b3005 := ("10" = r2984(0 to 1));
                                      goto_L3007 := b3005;
                                      if (NOT goto_L3007) then
                                        goto_L3013 := (NOT b3005);
                                        null; -- label L3013
                                        -- alt exit (no match)
                                        -- final pat
                                        -- got s@FA in r2980
                                        -- got vD'@F9 in r2978
                                        r3017 := rewire_setR3_1349(r2980,r2978);
                                        statevar0 := r3017;
                                        null;
                                        goto_L2986 := true;
                                      end if;
                                      goto_L2986 := goto_L2986;
                                      if (NOT goto_L2986) then
                                        null; -- label L3007
                                        -- got s@FA in r2980
                                        -- got vD'@F9 in r2978
                                        r3009 := rewire_setR2_1306(r2980,r2978);
                                        statevar0 := r3009;
                                        null;
                                        goto_L2986 := true;
                                      end if;
                                      goto_L2986 := goto_L2986;
                                    end if;
                                    goto_L2986 := goto_L2986;
                                    if (NOT goto_L2986) then
                                      null; -- label L2998
                                      -- got s@FA in r2980
                                      -- got vD'@F9 in r2978
                                      r3000 := rewire_setR1_1262(r2980,r2978);
                                      statevar0 := r3000;
                                      null;
                                      goto_L2986 := true;
                                    end if;
                                    goto_L2986 := goto_L2986;
                                  end if;
                                  goto_L2986 := goto_L2986;
                                  if (NOT goto_L2986) then
                                    null; -- label L2989
                                    -- got s@FA in r2980
                                    -- got vD'@F9 in r2978
                                    r2991 := rewire_setR0_1218(r2980,r2978);
                                    statevar0 := r2991;
                                    null;
                                    goto_L2986 := true;
                                  end if;
                                  goto_L2986 := goto_L2986;
                                  null; -- label L2986
                                  -- end case
                                  r3021 := statevar0;
                                  -- got s@FC in r3021
                                  r3024 := "0";
                                  r3026 := rewire_setCFlag_5(r3021,r3024);
                                  statevar0 := r3026;
                                  r3029 := statevar0;
                                  -- got s@FE in r3029
                                  -- got vD'@F9 in r2978
                                  r3033 := zeroW8;
                                  r3035 := eqW8(r2978,r3033);
                                  r3037 := rewire_setZFlag_48(r3029,r3035);
                                  statevar0 := r3037;
                                  r3040 := statevar0;
                                  -- got s@FG in r3040
                                  r3043 := rewire_outputs_144(r3040);
                                  -- got o@FH in r3043
                                  nextout := r3043;
                                  state := STATE3048;
                                  goto_L5439 := true;
                                end if;
                                goto_L5439 := goto_L5439;
                              end if;
                              goto_L5439 := goto_L5439;
                              if (NOT goto_L5439) then
                                null; -- label L2723
                                r2722 := statevar0;
                                -- got b0@EE in r2696
                                -- got b1@EF in r2698
                                r2726 := rewire_mkReg_883(r2696,r2698);
                                b2730 := ("00" = r2726(0 to 1));
                                goto_L2732 := b2730;
                                if (NOT goto_L2732) then
                                  goto_L2736 := (NOT b2730);
                                  null; -- label L2736
                                  -- alt exit (no match)
                                  b2737 := ("01" = r2726(0 to 1));
                                  goto_L2739 := b2737;
                                  if (NOT goto_L2739) then
                                    goto_L2743 := (NOT b2737);
                                    null; -- label L2743
                                    -- alt exit (no match)
                                    b2744 := ("10" = r2726(0 to 1));
                                    goto_L2746 := b2744;
                                    if (NOT goto_L2746) then
                                      goto_L2750 := (NOT b2744);
                                      null; -- label L2750
                                      -- alt exit (no match)
                                      -- final pat
                                      -- got s@EI in r2722
                                      r2753 := rewire_r3_1046(r2722);
                                      r2728 := r2753;
                                      goto_L2729 := true;
                                    end if;
                                    goto_L2729 := goto_L2729;
                                    if (NOT goto_L2729) then
                                      null; -- label L2746
                                      -- got s@EI in r2722
                                      r2747 := rewire_r2_1008(r2722);
                                      r2728 := r2747;
                                      goto_L2729 := true;
                                    end if;
                                    goto_L2729 := goto_L2729;
                                  end if;
                                  goto_L2729 := goto_L2729;
                                  if (NOT goto_L2729) then
                                    null; -- label L2739
                                    -- got s@EI in r2722
                                    r2740 := rewire_r1_969(r2722);
                                    r2728 := r2740;
                                    goto_L2729 := true;
                                  end if;
                                  goto_L2729 := goto_L2729;
                                end if;
                                goto_L2729 := goto_L2729;
                                if (NOT goto_L2729) then
                                  null; -- label L2732
                                  -- got s@EI in r2722
                                  r2733 := rewire_r0_930(r2722);
                                  r2728 := r2733;
                                  goto_L2729 := true;
                                end if;
                                goto_L2729 := goto_L2729;
                                null; -- label L2729
                                -- end case
                                r2756 := statevar0;
                                -- got c0@EG in r2700
                                -- got c1@EH in r2702
                                r2760 := rewire_mkReg_883(r2700,r2702);
                                b2764 := ("00" = r2760(0 to 1));
                                goto_L2766 := b2764;
                                if (NOT goto_L2766) then
                                  goto_L2770 := (NOT b2764);
                                  null; -- label L2770
                                  -- alt exit (no match)
                                  b2771 := ("01" = r2760(0 to 1));
                                  goto_L2773 := b2771;
                                  if (NOT goto_L2773) then
                                    goto_L2777 := (NOT b2771);
                                    null; -- label L2777
                                    -- alt exit (no match)
                                    b2778 := ("10" = r2760(0 to 1));
                                    goto_L2780 := b2778;
                                    if (NOT goto_L2780) then
                                      goto_L2784 := (NOT b2778);
                                      null; -- label L2784
                                      -- alt exit (no match)
                                      -- final pat
                                      -- got s@EK in r2756
                                      r2787 := rewire_r3_1046(r2756);
                                      r2762 := r2787;
                                      goto_L2763 := true;
                                    end if;
                                    goto_L2763 := goto_L2763;
                                    if (NOT goto_L2763) then
                                      null; -- label L2780
                                      -- got s@EK in r2756
                                      r2781 := rewire_r2_1008(r2756);
                                      r2762 := r2781;
                                      goto_L2763 := true;
                                    end if;
                                    goto_L2763 := goto_L2763;
                                  end if;
                                  goto_L2763 := goto_L2763;
                                  if (NOT goto_L2763) then
                                    null; -- label L2773
                                    -- got s@EK in r2756
                                    r2774 := rewire_r1_969(r2756);
                                    r2762 := r2774;
                                    goto_L2763 := true;
                                  end if;
                                  goto_L2763 := goto_L2763;
                                end if;
                                goto_L2763 := goto_L2763;
                                if (NOT goto_L2763) then
                                  null; -- label L2766
                                  -- got s@EK in r2756
                                  r2767 := rewire_r0_930(r2756);
                                  r2762 := r2767;
                                  goto_L2763 := true;
                                end if;
                                goto_L2763 := goto_L2763;
                                null; -- label L2763
                                -- end case
                                -- got vD@EJ in r2728
                                -- got vS@EL in r2762
                                r2792 := orW8(r2728,r2762);
                                r2794 := statevar0;
                                -- got b0@EE in r2696
                                -- got b1@EF in r2698
                                r2798 := rewire_mkReg_883(r2696,r2698);
                                b2801 := ("00" = r2798(0 to 1));
                                goto_L2803 := b2801;
                                if (NOT goto_L2803) then
                                  goto_L2809 := (NOT b2801);
                                  null; -- label L2809
                                  -- alt exit (no match)
                                  b2810 := ("01" = r2798(0 to 1));
                                  goto_L2812 := b2810;
                                  if (NOT goto_L2812) then
                                    goto_L2818 := (NOT b2810);
                                    null; -- label L2818
                                    -- alt exit (no match)
                                    b2819 := ("10" = r2798(0 to 1));
                                    goto_L2821 := b2819;
                                    if (NOT goto_L2821) then
                                      goto_L2827 := (NOT b2819);
                                      null; -- label L2827
                                      -- alt exit (no match)
                                      -- final pat
                                      -- got s@EN in r2794
                                      -- got vD'@EM in r2792
                                      r2831 := rewire_setR3_1349(r2794,r2792);
                                      statevar0 := r2831;
                                      null;
                                      goto_L2800 := true;
                                    end if;
                                    goto_L2800 := goto_L2800;
                                    if (NOT goto_L2800) then
                                      null; -- label L2821
                                      -- got s@EN in r2794
                                      -- got vD'@EM in r2792
                                      r2823 := rewire_setR2_1306(r2794,r2792);
                                      statevar0 := r2823;
                                      null;
                                      goto_L2800 := true;
                                    end if;
                                    goto_L2800 := goto_L2800;
                                  end if;
                                  goto_L2800 := goto_L2800;
                                  if (NOT goto_L2800) then
                                    null; -- label L2812
                                    -- got s@EN in r2794
                                    -- got vD'@EM in r2792
                                    r2814 := rewire_setR1_1262(r2794,r2792);
                                    statevar0 := r2814;
                                    null;
                                    goto_L2800 := true;
                                  end if;
                                  goto_L2800 := goto_L2800;
                                end if;
                                goto_L2800 := goto_L2800;
                                if (NOT goto_L2800) then
                                  null; -- label L2803
                                  -- got s@EN in r2794
                                  -- got vD'@EM in r2792
                                  r2805 := rewire_setR0_1218(r2794,r2792);
                                  statevar0 := r2805;
                                  null;
                                  goto_L2800 := true;
                                end if;
                                goto_L2800 := goto_L2800;
                                null; -- label L2800
                                -- end case
                                r2835 := statevar0;
                                -- got s@EP in r2835
                                r2838 := "0";
                                r2840 := rewire_setCFlag_5(r2835,r2838);
                                statevar0 := r2840;
                                r2843 := statevar0;
                                -- got s@ER in r2843
                                -- got vD'@EM in r2792
                                r2847 := zeroW8;
                                r2849 := eqW8(r2792,r2847);
                                r2851 := rewire_setZFlag_48(r2843,r2849);
                                statevar0 := r2851;
                                r2854 := statevar0;
                                -- got s@ET in r2854
                                r2857 := rewire_outputs_144(r2854);
                                -- got o@EU in r2857
                                nextout := r2857;
                                state := STATE2862;
                                goto_L5439 := true;
                              end if;
                              goto_L5439 := goto_L5439;
                            end if;
                            goto_L5439 := goto_L5439;
                            if (NOT goto_L5439) then
                              null; -- label L2594
                              r2593 := statevar0;
                              -- got c0@E4 in r2571
                              -- got c1@E5 in r2573
                              r2597 := rewire_mkReg_883(r2571,r2573);
                              b2601 := ("00" = r2597(0 to 1));
                              goto_L2603 := b2601;
                              if (NOT goto_L2603) then
                                goto_L2607 := (NOT b2601);
                                null; -- label L2607
                                -- alt exit (no match)
                                b2608 := ("01" = r2597(0 to 1));
                                goto_L2610 := b2608;
                                if (NOT goto_L2610) then
                                  goto_L2614 := (NOT b2608);
                                  null; -- label L2614
                                  -- alt exit (no match)
                                  b2615 := ("10" = r2597(0 to 1));
                                  goto_L2617 := b2615;
                                  if (NOT goto_L2617) then
                                    goto_L2621 := (NOT b2615);
                                    null; -- label L2621
                                    -- alt exit (no match)
                                    -- final pat
                                    -- got s@E6 in r2593
                                    r2624 := rewire_r3_1046(r2593);
                                    r2599 := r2624;
                                    goto_L2600 := true;
                                  end if;
                                  goto_L2600 := goto_L2600;
                                  if (NOT goto_L2600) then
                                    null; -- label L2617
                                    -- got s@E6 in r2593
                                    r2618 := rewire_r2_1008(r2593);
                                    r2599 := r2618;
                                    goto_L2600 := true;
                                  end if;
                                  goto_L2600 := goto_L2600;
                                end if;
                                goto_L2600 := goto_L2600;
                                if (NOT goto_L2600) then
                                  null; -- label L2610
                                  -- got s@E6 in r2593
                                  r2611 := rewire_r1_969(r2593);
                                  r2599 := r2611;
                                  goto_L2600 := true;
                                end if;
                                goto_L2600 := goto_L2600;
                              end if;
                              goto_L2600 := goto_L2600;
                              if (NOT goto_L2600) then
                                null; -- label L2603
                                -- got s@E6 in r2593
                                r2604 := rewire_r0_930(r2593);
                                r2599 := r2604;
                                goto_L2600 := true;
                              end if;
                              goto_L2600 := goto_L2600;
                              null; -- label L2600
                              -- end case
                              r2627 := statevar0;
                              -- got b0@E2 in r2567
                              -- got b1@E3 in r2569
                              r2631 := rewire_mkReg_883(r2567,r2569);
                              b2634 := ("00" = r2631(0 to 1));
                              goto_L2636 := b2634;
                              if (NOT goto_L2636) then
                                goto_L2642 := (NOT b2634);
                                null; -- label L2642
                                -- alt exit (no match)
                                b2643 := ("01" = r2631(0 to 1));
                                goto_L2645 := b2643;
                                if (NOT goto_L2645) then
                                  goto_L2651 := (NOT b2643);
                                  null; -- label L2651
                                  -- alt exit (no match)
                                  b2652 := ("10" = r2631(0 to 1));
                                  goto_L2654 := b2652;
                                  if (NOT goto_L2654) then
                                    goto_L2660 := (NOT b2652);
                                    null; -- label L2660
                                    -- alt exit (no match)
                                    -- final pat
                                    -- got s@E8 in r2627
                                    -- got v@E7 in r2599
                                    r2664 := rewire_setR3_1349(r2627,r2599);
                                    statevar0 := r2664;
                                    null;
                                    goto_L2633 := true;
                                  end if;
                                  goto_L2633 := goto_L2633;
                                  if (NOT goto_L2633) then
                                    null; -- label L2654
                                    -- got s@E8 in r2627
                                    -- got v@E7 in r2599
                                    r2656 := rewire_setR2_1306(r2627,r2599);
                                    statevar0 := r2656;
                                    null;
                                    goto_L2633 := true;
                                  end if;
                                  goto_L2633 := goto_L2633;
                                end if;
                                goto_L2633 := goto_L2633;
                                if (NOT goto_L2633) then
                                  null; -- label L2645
                                  -- got s@E8 in r2627
                                  -- got v@E7 in r2599
                                  r2647 := rewire_setR1_1262(r2627,r2599);
                                  statevar0 := r2647;
                                  null;
                                  goto_L2633 := true;
                                end if;
                                goto_L2633 := goto_L2633;
                              end if;
                              goto_L2633 := goto_L2633;
                              if (NOT goto_L2633) then
                                null; -- label L2636
                                -- got s@E8 in r2627
                                -- got v@E7 in r2599
                                r2638 := rewire_setR0_1218(r2627,r2599);
                                statevar0 := r2638;
                                null;
                                goto_L2633 := true;
                              end if;
                              goto_L2633 := goto_L2633;
                              null; -- label L2633
                              -- end case
                              r2668 := statevar0;
                              -- got s@EA in r2668
                              r2671 := rewire_outputs_144(r2668);
                              -- got o@EB in r2671
                              nextout := r2671;
                              state := STATE2676;
                              goto_L5439 := true;
                            end if;
                            goto_L5439 := goto_L5439;
                          end if;
                          goto_L5439 := goto_L5439;
                          if (NOT goto_L5439) then
                            null; -- label L2386
                            r2385 := statevar0;
                            -- got b0@DB in r2359
                            -- got b1@DC in r2361
                            r2389 := rewire_mkReg_883(r2359,r2361);
                            b2393 := ("00" = r2389(0 to 1));
                            goto_L2395 := b2393;
                            if (NOT goto_L2395) then
                              goto_L2399 := (NOT b2393);
                              null; -- label L2399
                              -- alt exit (no match)
                              b2400 := ("01" = r2389(0 to 1));
                              goto_L2402 := b2400;
                              if (NOT goto_L2402) then
                                goto_L2406 := (NOT b2400);
                                null; -- label L2406
                                -- alt exit (no match)
                                b2407 := ("10" = r2389(0 to 1));
                                goto_L2409 := b2407;
                                if (NOT goto_L2409) then
                                  goto_L2413 := (NOT b2407);
                                  null; -- label L2413
                                  -- alt exit (no match)
                                  -- final pat
                                  -- got s@DF in r2385
                                  r2416 := rewire_r3_1046(r2385);
                                  r2391 := r2416;
                                  goto_L2392 := true;
                                end if;
                                goto_L2392 := goto_L2392;
                                if (NOT goto_L2392) then
                                  null; -- label L2409
                                  -- got s@DF in r2385
                                  r2410 := rewire_r2_1008(r2385);
                                  r2391 := r2410;
                                  goto_L2392 := true;
                                end if;
                                goto_L2392 := goto_L2392;
                              end if;
                              goto_L2392 := goto_L2392;
                              if (NOT goto_L2392) then
                                null; -- label L2402
                                -- got s@DF in r2385
                                r2403 := rewire_r1_969(r2385);
                                r2391 := r2403;
                                goto_L2392 := true;
                              end if;
                              goto_L2392 := goto_L2392;
                            end if;
                            goto_L2392 := goto_L2392;
                            if (NOT goto_L2392) then
                              null; -- label L2395
                              -- got s@DF in r2385
                              r2396 := rewire_r0_930(r2385);
                              r2391 := r2396;
                              goto_L2392 := true;
                            end if;
                            goto_L2392 := goto_L2392;
                            null; -- label L2392
                            -- end case
                            r2419 := statevar0;
                            -- got c0@DD in r2363
                            -- got c1@DE in r2365
                            r2423 := rewire_mkReg_883(r2363,r2365);
                            b2427 := ("00" = r2423(0 to 1));
                            goto_L2429 := b2427;
                            if (NOT goto_L2429) then
                              goto_L2433 := (NOT b2427);
                              null; -- label L2433
                              -- alt exit (no match)
                              b2434 := ("01" = r2423(0 to 1));
                              goto_L2436 := b2434;
                              if (NOT goto_L2436) then
                                goto_L2440 := (NOT b2434);
                                null; -- label L2440
                                -- alt exit (no match)
                                b2441 := ("10" = r2423(0 to 1));
                                goto_L2443 := b2441;
                                if (NOT goto_L2443) then
                                  goto_L2447 := (NOT b2441);
                                  null; -- label L2447
                                  -- alt exit (no match)
                                  -- final pat
                                  -- got s@DH in r2419
                                  r2450 := rewire_r3_1046(r2419);
                                  r2425 := r2450;
                                  goto_L2426 := true;
                                end if;
                                goto_L2426 := goto_L2426;
                                if (NOT goto_L2426) then
                                  null; -- label L2443
                                  -- got s@DH in r2419
                                  r2444 := rewire_r2_1008(r2419);
                                  r2425 := r2444;
                                  goto_L2426 := true;
                                end if;
                                goto_L2426 := goto_L2426;
                              end if;
                              goto_L2426 := goto_L2426;
                              if (NOT goto_L2426) then
                                null; -- label L2436
                                -- got s@DH in r2419
                                r2437 := rewire_r1_969(r2419);
                                r2425 := r2437;
                                goto_L2426 := true;
                              end if;
                              goto_L2426 := goto_L2426;
                            end if;
                            goto_L2426 := goto_L2426;
                            if (NOT goto_L2426) then
                              null; -- label L2429
                              -- got s@DH in r2419
                              r2430 := rewire_r0_930(r2419);
                              r2425 := r2430;
                              goto_L2426 := true;
                            end if;
                            goto_L2426 := goto_L2426;
                            null; -- label L2426
                            -- end case
                            r2453 := statevar0;
                            -- got s@DJ in r2453
                            r2456 := rewire_cFlag_536(r2453);
                            -- got vD@DG in r2391
                            -- got vS@DI in r2425
                            -- got cin@DK in r2456
                            r2461 := minusCW8(r2391,r2425,r2456);
                            -- got p@DL in r2461
                            -- final pat
                            r2466 := r2461(0 to 0);
                            r2468 := r2461(1 to 8);
                            b2470 := true;
                            b2472 := true;
                            -- got x@DM in r2466
                            r2464 := r2466;
                            -- end case
                            -- got p@DL in r2461
                            -- final pat
                            r2480 := r2461(0 to 0);
                            r2482 := r2461(1 to 8);
                            b2484 := true;
                            b2486 := true;
                            -- got x@DO in r2482
                            r2478 := r2482;
                            -- end case
                            r2491 := statevar0;
                            -- got s@DQ in r2491
                            -- got cout@DN in r2464
                            r2495 := rewire_setCFlag_5(r2491,r2464);
                            statevar0 := r2495;
                            r2498 := statevar0;
                            -- got b0@DB in r2359
                            -- got b1@DC in r2361
                            r2502 := rewire_mkReg_883(r2359,r2361);
                            b2505 := ("00" = r2502(0 to 1));
                            goto_L2507 := b2505;
                            if (NOT goto_L2507) then
                              goto_L2513 := (NOT b2505);
                              null; -- label L2513
                              -- alt exit (no match)
                              b2514 := ("01" = r2502(0 to 1));
                              goto_L2516 := b2514;
                              if (NOT goto_L2516) then
                                goto_L2522 := (NOT b2514);
                                null; -- label L2522
                                -- alt exit (no match)
                                b2523 := ("10" = r2502(0 to 1));
                                goto_L2525 := b2523;
                                if (NOT goto_L2525) then
                                  goto_L2531 := (NOT b2523);
                                  null; -- label L2531
                                  -- alt exit (no match)
                                  -- final pat
                                  -- got s@DS in r2498
                                  -- got vD'@DP in r2478
                                  r2535 := rewire_setR3_1349(r2498,r2478);
                                  statevar0 := r2535;
                                  null;
                                  goto_L2504 := true;
                                end if;
                                goto_L2504 := goto_L2504;
                                if (NOT goto_L2504) then
                                  null; -- label L2525
                                  -- got s@DS in r2498
                                  -- got vD'@DP in r2478
                                  r2527 := rewire_setR2_1306(r2498,r2478);
                                  statevar0 := r2527;
                                  null;
                                  goto_L2504 := true;
                                end if;
                                goto_L2504 := goto_L2504;
                              end if;
                              goto_L2504 := goto_L2504;
                              if (NOT goto_L2504) then
                                null; -- label L2516
                                -- got s@DS in r2498
                                -- got vD'@DP in r2478
                                r2518 := rewire_setR1_1262(r2498,r2478);
                                statevar0 := r2518;
                                null;
                                goto_L2504 := true;
                              end if;
                              goto_L2504 := goto_L2504;
                            end if;
                            goto_L2504 := goto_L2504;
                            if (NOT goto_L2504) then
                              null; -- label L2507
                              -- got s@DS in r2498
                              -- got vD'@DP in r2478
                              r2509 := rewire_setR0_1218(r2498,r2478);
                              statevar0 := r2509;
                              null;
                              goto_L2504 := true;
                            end if;
                            goto_L2504 := goto_L2504;
                            null; -- label L2504
                            -- end case
                            r2539 := statevar0;
                            -- got s@DU in r2539
                            r2542 := rewire_outputs_144(r2539);
                            -- got o@DV in r2542
                            nextout := r2542;
                            state := STATE2547;
                            goto_L5439 := true;
                          end if;
                          goto_L5439 := goto_L5439;
                        end if;
                        goto_L5439 := goto_L5439;
                        if (NOT goto_L5439) then
                          null; -- label L2182
                          r2181 := statevar0;
                          -- got b0@CM in r2155
                          -- got b1@CN in r2157
                          r2185 := rewire_mkReg_883(r2155,r2157);
                          b2189 := ("00" = r2185(0 to 1));
                          goto_L2191 := b2189;
                          if (NOT goto_L2191) then
                            goto_L2195 := (NOT b2189);
                            null; -- label L2195
                            -- alt exit (no match)
                            b2196 := ("01" = r2185(0 to 1));
                            goto_L2198 := b2196;
                            if (NOT goto_L2198) then
                              goto_L2202 := (NOT b2196);
                              null; -- label L2202
                              -- alt exit (no match)
                              b2203 := ("10" = r2185(0 to 1));
                              goto_L2205 := b2203;
                              if (NOT goto_L2205) then
                                goto_L2209 := (NOT b2203);
                                null; -- label L2209
                                -- alt exit (no match)
                                -- final pat
                                -- got s@CQ in r2181
                                r2212 := rewire_r3_1046(r2181);
                                r2187 := r2212;
                                goto_L2188 := true;
                              end if;
                              goto_L2188 := goto_L2188;
                              if (NOT goto_L2188) then
                                null; -- label L2205
                                -- got s@CQ in r2181
                                r2206 := rewire_r2_1008(r2181);
                                r2187 := r2206;
                                goto_L2188 := true;
                              end if;
                              goto_L2188 := goto_L2188;
                            end if;
                            goto_L2188 := goto_L2188;
                            if (NOT goto_L2188) then
                              null; -- label L2198
                              -- got s@CQ in r2181
                              r2199 := rewire_r1_969(r2181);
                              r2187 := r2199;
                              goto_L2188 := true;
                            end if;
                            goto_L2188 := goto_L2188;
                          end if;
                          goto_L2188 := goto_L2188;
                          if (NOT goto_L2188) then
                            null; -- label L2191
                            -- got s@CQ in r2181
                            r2192 := rewire_r0_930(r2181);
                            r2187 := r2192;
                            goto_L2188 := true;
                          end if;
                          goto_L2188 := goto_L2188;
                          null; -- label L2188
                          -- end case
                          r2215 := statevar0;
                          -- got c0@CO in r2159
                          -- got c1@CP in r2161
                          r2219 := rewire_mkReg_883(r2159,r2161);
                          b2223 := ("00" = r2219(0 to 1));
                          goto_L2225 := b2223;
                          if (NOT goto_L2225) then
                            goto_L2229 := (NOT b2223);
                            null; -- label L2229
                            -- alt exit (no match)
                            b2230 := ("01" = r2219(0 to 1));
                            goto_L2232 := b2230;
                            if (NOT goto_L2232) then
                              goto_L2236 := (NOT b2230);
                              null; -- label L2236
                              -- alt exit (no match)
                              b2237 := ("10" = r2219(0 to 1));
                              goto_L2239 := b2237;
                              if (NOT goto_L2239) then
                                goto_L2243 := (NOT b2237);
                                null; -- label L2243
                                -- alt exit (no match)
                                -- final pat
                                -- got s@CS in r2215
                                r2246 := rewire_r3_1046(r2215);
                                r2221 := r2246;
                                goto_L2222 := true;
                              end if;
                              goto_L2222 := goto_L2222;
                              if (NOT goto_L2222) then
                                null; -- label L2239
                                -- got s@CS in r2215
                                r2240 := rewire_r2_1008(r2215);
                                r2221 := r2240;
                                goto_L2222 := true;
                              end if;
                              goto_L2222 := goto_L2222;
                            end if;
                            goto_L2222 := goto_L2222;
                            if (NOT goto_L2222) then
                              null; -- label L2232
                              -- got s@CS in r2215
                              r2233 := rewire_r1_969(r2215);
                              r2221 := r2233;
                              goto_L2222 := true;
                            end if;
                            goto_L2222 := goto_L2222;
                          end if;
                          goto_L2222 := goto_L2222;
                          if (NOT goto_L2222) then
                            null; -- label L2225
                            -- got s@CS in r2215
                            r2226 := rewire_r0_930(r2215);
                            r2221 := r2226;
                            goto_L2222 := true;
                          end if;
                          goto_L2222 := goto_L2222;
                          null; -- label L2222
                          -- end case
                          -- got vD@CR in r2187
                          -- got vS@CT in r2221
                          r2251 := "0";
                          r2253 := minusCW8(r2187,r2221,r2251);
                          -- got p@CU in r2253
                          -- final pat
                          r2258 := r2253(0 to 0);
                          r2260 := r2253(1 to 8);
                          b2262 := true;
                          b2264 := true;
                          -- got x@CV in r2258
                          r2256 := r2258;
                          -- end case
                          -- got p@CU in r2253
                          -- final pat
                          r2272 := r2253(0 to 0);
                          r2274 := r2253(1 to 8);
                          b2276 := true;
                          b2278 := true;
                          -- got x@D1 in r2274
                          r2270 := r2274;
                          -- end case
                          r2283 := statevar0;
                          -- got s@D3 in r2283
                          -- got cout@D0 in r2256
                          r2287 := rewire_setCFlag_5(r2283,r2256);
                          statevar0 := r2287;
                          r2290 := statevar0;
                          -- got b0@CM in r2155
                          -- got b1@CN in r2157
                          r2294 := rewire_mkReg_883(r2155,r2157);
                          b2297 := ("00" = r2294(0 to 1));
                          goto_L2299 := b2297;
                          if (NOT goto_L2299) then
                            goto_L2305 := (NOT b2297);
                            null; -- label L2305
                            -- alt exit (no match)
                            b2306 := ("01" = r2294(0 to 1));
                            goto_L2308 := b2306;
                            if (NOT goto_L2308) then
                              goto_L2314 := (NOT b2306);
                              null; -- label L2314
                              -- alt exit (no match)
                              b2315 := ("10" = r2294(0 to 1));
                              goto_L2317 := b2315;
                              if (NOT goto_L2317) then
                                goto_L2323 := (NOT b2315);
                                null; -- label L2323
                                -- alt exit (no match)
                                -- final pat
                                -- got s@D5 in r2290
                                -- got vD'@D2 in r2270
                                r2327 := rewire_setR3_1349(r2290,r2270);
                                statevar0 := r2327;
                                null;
                                goto_L2296 := true;
                              end if;
                              goto_L2296 := goto_L2296;
                              if (NOT goto_L2296) then
                                null; -- label L2317
                                -- got s@D5 in r2290
                                -- got vD'@D2 in r2270
                                r2319 := rewire_setR2_1306(r2290,r2270);
                                statevar0 := r2319;
                                null;
                                goto_L2296 := true;
                              end if;
                              goto_L2296 := goto_L2296;
                            end if;
                            goto_L2296 := goto_L2296;
                            if (NOT goto_L2296) then
                              null; -- label L2308
                              -- got s@D5 in r2290
                              -- got vD'@D2 in r2270
                              r2310 := rewire_setR1_1262(r2290,r2270);
                              statevar0 := r2310;
                              null;
                              goto_L2296 := true;
                            end if;
                            goto_L2296 := goto_L2296;
                          end if;
                          goto_L2296 := goto_L2296;
                          if (NOT goto_L2296) then
                            null; -- label L2299
                            -- got s@D5 in r2290
                            -- got vD'@D2 in r2270
                            r2301 := rewire_setR0_1218(r2290,r2270);
                            statevar0 := r2301;
                            null;
                            goto_L2296 := true;
                          end if;
                          goto_L2296 := goto_L2296;
                          null; -- label L2296
                          -- end case
                          r2331 := statevar0;
                          -- got s@D7 in r2331
                          r2334 := rewire_outputs_144(r2331);
                          -- got o@D8 in r2334
                          nextout := r2334;
                          state := STATE2339;
                          goto_L5439 := true;
                        end if;
                        goto_L5439 := goto_L5439;
                      end if;
                      goto_L5439 := goto_L5439;
                      if (NOT goto_L5439) then
                        null; -- label L1974
                        r1973 := statevar0;
                        -- got b0@BV in r1947
                        -- got b1@C0 in r1949
                        r1977 := rewire_mkReg_883(r1947,r1949);
                        b1981 := ("00" = r1977(0 to 1));
                        goto_L1983 := b1981;
                        if (NOT goto_L1983) then
                          goto_L1987 := (NOT b1981);
                          null; -- label L1987
                          -- alt exit (no match)
                          b1988 := ("01" = r1977(0 to 1));
                          goto_L1990 := b1988;
                          if (NOT goto_L1990) then
                            goto_L1994 := (NOT b1988);
                            null; -- label L1994
                            -- alt exit (no match)
                            b1995 := ("10" = r1977(0 to 1));
                            goto_L1997 := b1995;
                            if (NOT goto_L1997) then
                              goto_L2001 := (NOT b1995);
                              null; -- label L2001
                              -- alt exit (no match)
                              -- final pat
                              -- got s@C3 in r1973
                              r2004 := rewire_r3_1046(r1973);
                              r1979 := r2004;
                              goto_L1980 := true;
                            end if;
                            goto_L1980 := goto_L1980;
                            if (NOT goto_L1980) then
                              null; -- label L1997
                              -- got s@C3 in r1973
                              r1998 := rewire_r2_1008(r1973);
                              r1979 := r1998;
                              goto_L1980 := true;
                            end if;
                            goto_L1980 := goto_L1980;
                          end if;
                          goto_L1980 := goto_L1980;
                          if (NOT goto_L1980) then
                            null; -- label L1990
                            -- got s@C3 in r1973
                            r1991 := rewire_r1_969(r1973);
                            r1979 := r1991;
                            goto_L1980 := true;
                          end if;
                          goto_L1980 := goto_L1980;
                        end if;
                        goto_L1980 := goto_L1980;
                        if (NOT goto_L1980) then
                          null; -- label L1983
                          -- got s@C3 in r1973
                          r1984 := rewire_r0_930(r1973);
                          r1979 := r1984;
                          goto_L1980 := true;
                        end if;
                        goto_L1980 := goto_L1980;
                        null; -- label L1980
                        -- end case
                        r2007 := statevar0;
                        -- got c0@C1 in r1951
                        -- got c1@C2 in r1953
                        r2011 := rewire_mkReg_883(r1951,r1953);
                        b2015 := ("00" = r2011(0 to 1));
                        goto_L2017 := b2015;
                        if (NOT goto_L2017) then
                          goto_L2021 := (NOT b2015);
                          null; -- label L2021
                          -- alt exit (no match)
                          b2022 := ("01" = r2011(0 to 1));
                          goto_L2024 := b2022;
                          if (NOT goto_L2024) then
                            goto_L2028 := (NOT b2022);
                            null; -- label L2028
                            -- alt exit (no match)
                            b2029 := ("10" = r2011(0 to 1));
                            goto_L2031 := b2029;
                            if (NOT goto_L2031) then
                              goto_L2035 := (NOT b2029);
                              null; -- label L2035
                              -- alt exit (no match)
                              -- final pat
                              -- got s@C5 in r2007
                              r2038 := rewire_r3_1046(r2007);
                              r2013 := r2038;
                              goto_L2014 := true;
                            end if;
                            goto_L2014 := goto_L2014;
                            if (NOT goto_L2014) then
                              null; -- label L2031
                              -- got s@C5 in r2007
                              r2032 := rewire_r2_1008(r2007);
                              r2013 := r2032;
                              goto_L2014 := true;
                            end if;
                            goto_L2014 := goto_L2014;
                          end if;
                          goto_L2014 := goto_L2014;
                          if (NOT goto_L2014) then
                            null; -- label L2024
                            -- got s@C5 in r2007
                            r2025 := rewire_r1_969(r2007);
                            r2013 := r2025;
                            goto_L2014 := true;
                          end if;
                          goto_L2014 := goto_L2014;
                        end if;
                        goto_L2014 := goto_L2014;
                        if (NOT goto_L2014) then
                          null; -- label L2017
                          -- got s@C5 in r2007
                          r2018 := rewire_r0_930(r2007);
                          r2013 := r2018;
                          goto_L2014 := true;
                        end if;
                        goto_L2014 := goto_L2014;
                        null; -- label L2014
                        -- end case
                        r2041 := statevar0;
                        -- got s@C7 in r2041
                        r2044 := rewire_cFlag_536(r2041);
                        -- got vD@C4 in r1979
                        -- got vS@C6 in r2013
                        -- got cin@C8 in r2044
                        r2049 := plusCW8(r1979,r2013,r2044);
                        -- got p@C9 in r2049
                        -- final pat
                        r2054 := r2049(0 to 0);
                        r2056 := r2049(1 to 8);
                        b2058 := true;
                        b2060 := true;
                        -- got x@CA in r2054
                        r2052 := r2054;
                        -- end case
                        -- got p@C9 in r2049
                        -- final pat
                        r2068 := r2049(0 to 0);
                        r2070 := r2049(1 to 8);
                        b2072 := true;
                        b2074 := true;
                        -- got x@CC in r2070
                        r2066 := r2070;
                        -- end case
                        r2079 := statevar0;
                        -- got s@CE in r2079
                        -- got cout@CB in r2052
                        r2083 := rewire_setCFlag_5(r2079,r2052);
                        statevar0 := r2083;
                        r2086 := statevar0;
                        -- got b0@BV in r1947
                        -- got b1@C0 in r1949
                        r2090 := rewire_mkReg_883(r1947,r1949);
                        b2093 := ("00" = r2090(0 to 1));
                        goto_L2095 := b2093;
                        if (NOT goto_L2095) then
                          goto_L2101 := (NOT b2093);
                          null; -- label L2101
                          -- alt exit (no match)
                          b2102 := ("01" = r2090(0 to 1));
                          goto_L2104 := b2102;
                          if (NOT goto_L2104) then
                            goto_L2110 := (NOT b2102);
                            null; -- label L2110
                            -- alt exit (no match)
                            b2111 := ("10" = r2090(0 to 1));
                            goto_L2113 := b2111;
                            if (NOT goto_L2113) then
                              goto_L2119 := (NOT b2111);
                              null; -- label L2119
                              -- alt exit (no match)
                              -- final pat
                              -- got s@CG in r2086
                              -- got vD'@CD in r2066
                              r2123 := rewire_setR3_1349(r2086,r2066);
                              statevar0 := r2123;
                              null;
                              goto_L2092 := true;
                            end if;
                            goto_L2092 := goto_L2092;
                            if (NOT goto_L2092) then
                              null; -- label L2113
                              -- got s@CG in r2086
                              -- got vD'@CD in r2066
                              r2115 := rewire_setR2_1306(r2086,r2066);
                              statevar0 := r2115;
                              null;
                              goto_L2092 := true;
                            end if;
                            goto_L2092 := goto_L2092;
                          end if;
                          goto_L2092 := goto_L2092;
                          if (NOT goto_L2092) then
                            null; -- label L2104
                            -- got s@CG in r2086
                            -- got vD'@CD in r2066
                            r2106 := rewire_setR1_1262(r2086,r2066);
                            statevar0 := r2106;
                            null;
                            goto_L2092 := true;
                          end if;
                          goto_L2092 := goto_L2092;
                        end if;
                        goto_L2092 := goto_L2092;
                        if (NOT goto_L2092) then
                          null; -- label L2095
                          -- got s@CG in r2086
                          -- got vD'@CD in r2066
                          r2097 := rewire_setR0_1218(r2086,r2066);
                          statevar0 := r2097;
                          null;
                          goto_L2092 := true;
                        end if;
                        goto_L2092 := goto_L2092;
                        null; -- label L2092
                        -- end case
                        r2127 := statevar0;
                        -- got s@CI in r2127
                        r2130 := rewire_outputs_144(r2127);
                        -- got o@CJ in r2130
                        nextout := r2130;
                        state := STATE2135;
                        goto_L5439 := true;
                      end if;
                      goto_L5439 := goto_L5439;
                    end if;
                    goto_L5439 := goto_L5439;
                    if (NOT goto_L5439) then
                      null; -- label L1770
                      r1769 := statevar0;
                      -- got b0@BA in r1743
                      -- got b1@BB in r1745
                      r1773 := rewire_mkReg_883(r1743,r1745);
                      b1777 := ("00" = r1773(0 to 1));
                      goto_L1779 := b1777;
                      if (NOT goto_L1779) then
                        goto_L1783 := (NOT b1777);
                        null; -- label L1783
                        -- alt exit (no match)
                        b1784 := ("01" = r1773(0 to 1));
                        goto_L1786 := b1784;
                        if (NOT goto_L1786) then
                          goto_L1790 := (NOT b1784);
                          null; -- label L1790
                          -- alt exit (no match)
                          b1791 := ("10" = r1773(0 to 1));
                          goto_L1793 := b1791;
                          if (NOT goto_L1793) then
                            goto_L1797 := (NOT b1791);
                            null; -- label L1797
                            -- alt exit (no match)
                            -- final pat
                            -- got s@BE in r1769
                            r1800 := rewire_r3_1046(r1769);
                            r1775 := r1800;
                            goto_L1776 := true;
                          end if;
                          goto_L1776 := goto_L1776;
                          if (NOT goto_L1776) then
                            null; -- label L1793
                            -- got s@BE in r1769
                            r1794 := rewire_r2_1008(r1769);
                            r1775 := r1794;
                            goto_L1776 := true;
                          end if;
                          goto_L1776 := goto_L1776;
                        end if;
                        goto_L1776 := goto_L1776;
                        if (NOT goto_L1776) then
                          null; -- label L1786
                          -- got s@BE in r1769
                          r1787 := rewire_r1_969(r1769);
                          r1775 := r1787;
                          goto_L1776 := true;
                        end if;
                        goto_L1776 := goto_L1776;
                      end if;
                      goto_L1776 := goto_L1776;
                      if (NOT goto_L1776) then
                        null; -- label L1779
                        -- got s@BE in r1769
                        r1780 := rewire_r0_930(r1769);
                        r1775 := r1780;
                        goto_L1776 := true;
                      end if;
                      goto_L1776 := goto_L1776;
                      null; -- label L1776
                      -- end case
                      r1803 := statevar0;
                      -- got c0@BC in r1747
                      -- got c1@BD in r1749
                      r1807 := rewire_mkReg_883(r1747,r1749);
                      b1811 := ("00" = r1807(0 to 1));
                      goto_L1813 := b1811;
                      if (NOT goto_L1813) then
                        goto_L1817 := (NOT b1811);
                        null; -- label L1817
                        -- alt exit (no match)
                        b1818 := ("01" = r1807(0 to 1));
                        goto_L1820 := b1818;
                        if (NOT goto_L1820) then
                          goto_L1824 := (NOT b1818);
                          null; -- label L1824
                          -- alt exit (no match)
                          b1825 := ("10" = r1807(0 to 1));
                          goto_L1827 := b1825;
                          if (NOT goto_L1827) then
                            goto_L1831 := (NOT b1825);
                            null; -- label L1831
                            -- alt exit (no match)
                            -- final pat
                            -- got s@BG in r1803
                            r1834 := rewire_r3_1046(r1803);
                            r1809 := r1834;
                            goto_L1810 := true;
                          end if;
                          goto_L1810 := goto_L1810;
                          if (NOT goto_L1810) then
                            null; -- label L1827
                            -- got s@BG in r1803
                            r1828 := rewire_r2_1008(r1803);
                            r1809 := r1828;
                            goto_L1810 := true;
                          end if;
                          goto_L1810 := goto_L1810;
                        end if;
                        goto_L1810 := goto_L1810;
                        if (NOT goto_L1810) then
                          null; -- label L1820
                          -- got s@BG in r1803
                          r1821 := rewire_r1_969(r1803);
                          r1809 := r1821;
                          goto_L1810 := true;
                        end if;
                        goto_L1810 := goto_L1810;
                      end if;
                      goto_L1810 := goto_L1810;
                      if (NOT goto_L1810) then
                        null; -- label L1813
                        -- got s@BG in r1803
                        r1814 := rewire_r0_930(r1803);
                        r1809 := r1814;
                        goto_L1810 := true;
                      end if;
                      goto_L1810 := goto_L1810;
                      null; -- label L1810
                      -- end case
                      -- got vD@BF in r1775
                      -- got vS@BH in r1809
                      r1839 := "0";
                      r1841 := plusCW8(r1775,r1809,r1839);
                      -- got p@BI in r1841
                      -- final pat
                      r1846 := r1841(0 to 0);
                      r1848 := r1841(1 to 8);
                      b1850 := true;
                      b1852 := true;
                      -- got x@BJ in r1846
                      r1844 := r1846;
                      -- end case
                      -- got p@BI in r1841
                      -- final pat
                      r1860 := r1841(0 to 0);
                      r1862 := r1841(1 to 8);
                      b1864 := true;
                      b1866 := true;
                      -- got x@BL in r1862
                      r1858 := r1862;
                      -- end case
                      r1871 := statevar0;
                      -- got s@BN in r1871
                      -- got cout@BK in r1844
                      r1875 := rewire_setCFlag_5(r1871,r1844);
                      statevar0 := r1875;
                      r1878 := statevar0;
                      -- got b0@BA in r1743
                      -- got b1@BB in r1745
                      r1882 := rewire_mkReg_883(r1743,r1745);
                      b1885 := ("00" = r1882(0 to 1));
                      goto_L1887 := b1885;
                      if (NOT goto_L1887) then
                        goto_L1893 := (NOT b1885);
                        null; -- label L1893
                        -- alt exit (no match)
                        b1894 := ("01" = r1882(0 to 1));
                        goto_L1896 := b1894;
                        if (NOT goto_L1896) then
                          goto_L1902 := (NOT b1894);
                          null; -- label L1902
                          -- alt exit (no match)
                          b1903 := ("10" = r1882(0 to 1));
                          goto_L1905 := b1903;
                          if (NOT goto_L1905) then
                            goto_L1911 := (NOT b1903);
                            null; -- label L1911
                            -- alt exit (no match)
                            -- final pat
                            -- got s@BP in r1878
                            -- got vD'@BM in r1858
                            r1915 := rewire_setR3_1349(r1878,r1858);
                            statevar0 := r1915;
                            null;
                            goto_L1884 := true;
                          end if;
                          goto_L1884 := goto_L1884;
                          if (NOT goto_L1884) then
                            null; -- label L1905
                            -- got s@BP in r1878
                            -- got vD'@BM in r1858
                            r1907 := rewire_setR2_1306(r1878,r1858);
                            statevar0 := r1907;
                            null;
                            goto_L1884 := true;
                          end if;
                          goto_L1884 := goto_L1884;
                        end if;
                        goto_L1884 := goto_L1884;
                        if (NOT goto_L1884) then
                          null; -- label L1896
                          -- got s@BP in r1878
                          -- got vD'@BM in r1858
                          r1898 := rewire_setR1_1262(r1878,r1858);
                          statevar0 := r1898;
                          null;
                          goto_L1884 := true;
                        end if;
                        goto_L1884 := goto_L1884;
                      end if;
                      goto_L1884 := goto_L1884;
                      if (NOT goto_L1884) then
                        null; -- label L1887
                        -- got s@BP in r1878
                        -- got vD'@BM in r1858
                        r1889 := rewire_setR0_1218(r1878,r1858);
                        statevar0 := r1889;
                        null;
                        goto_L1884 := true;
                      end if;
                      goto_L1884 := goto_L1884;
                      null; -- label L1884
                      -- end case
                      r1919 := statevar0;
                      -- got s@BR in r1919
                      r1922 := rewire_outputs_144(r1919);
                      -- got o@BS in r1922
                      nextout := r1922;
                      state := STATE1927;
                      goto_L5439 := true;
                    end if;
                    goto_L5439 := goto_L5439;
                  end if;
                  goto_L5439 := goto_L5439;
                  if (NOT goto_L5439) then
                    null; -- label L1602
                    r1601 := statevar0;
                    -- got c0@AK in r1579
                    -- got c1@AL in r1581
                    r1605 := rewire_mkReg_883(r1579,r1581);
                    b1609 := ("00" = r1605(0 to 1));
                    goto_L1611 := b1609;
                    if (NOT goto_L1611) then
                      goto_L1615 := (NOT b1609);
                      null; -- label L1615
                      -- alt exit (no match)
                      b1616 := ("01" = r1605(0 to 1));
                      goto_L1618 := b1616;
                      if (NOT goto_L1618) then
                        goto_L1622 := (NOT b1616);
                        null; -- label L1622
                        -- alt exit (no match)
                        b1623 := ("10" = r1605(0 to 1));
                        goto_L1625 := b1623;
                        if (NOT goto_L1625) then
                          goto_L1629 := (NOT b1623);
                          null; -- label L1629
                          -- alt exit (no match)
                          -- final pat
                          -- got s@AM in r1601
                          r1632 := rewire_r3_1046(r1601);
                          r1607 := r1632;
                          goto_L1608 := true;
                        end if;
                        goto_L1608 := goto_L1608;
                        if (NOT goto_L1608) then
                          null; -- label L1625
                          -- got s@AM in r1601
                          r1626 := rewire_r2_1008(r1601);
                          r1607 := r1626;
                          goto_L1608 := true;
                        end if;
                        goto_L1608 := goto_L1608;
                      end if;
                      goto_L1608 := goto_L1608;
                      if (NOT goto_L1608) then
                        null; -- label L1618
                        -- got s@AM in r1601
                        r1619 := rewire_r1_969(r1601);
                        r1607 := r1619;
                        goto_L1608 := true;
                      end if;
                      goto_L1608 := goto_L1608;
                    end if;
                    goto_L1608 := goto_L1608;
                    if (NOT goto_L1608) then
                      null; -- label L1611
                      -- got s@AM in r1601
                      r1612 := rewire_r0_930(r1601);
                      r1607 := r1612;
                      goto_L1608 := true;
                    end if;
                    goto_L1608 := goto_L1608;
                    null; -- label L1608
                    -- end case
                    r1635 := statevar0;
                    -- got b0@AI in r1575
                    -- got b1@AJ in r1577
                    r1639 := rewire_mkReg_883(r1575,r1577);
                    b1643 := ("00" = r1639(0 to 1));
                    goto_L1645 := b1643;
                    if (NOT goto_L1645) then
                      goto_L1649 := (NOT b1643);
                      null; -- label L1649
                      -- alt exit (no match)
                      b1650 := ("01" = r1639(0 to 1));
                      goto_L1652 := b1650;
                      if (NOT goto_L1652) then
                        goto_L1656 := (NOT b1650);
                        null; -- label L1656
                        -- alt exit (no match)
                        b1657 := ("10" = r1639(0 to 1));
                        goto_L1659 := b1657;
                        if (NOT goto_L1659) then
                          goto_L1663 := (NOT b1657);
                          null; -- label L1663
                          -- alt exit (no match)
                          -- final pat
                          -- got s@AO in r1635
                          r1666 := rewire_r3_1046(r1635);
                          r1641 := r1666;
                          goto_L1642 := true;
                        end if;
                        goto_L1642 := goto_L1642;
                        if (NOT goto_L1642) then
                          null; -- label L1659
                          -- got s@AO in r1635
                          r1660 := rewire_r2_1008(r1635);
                          r1641 := r1660;
                          goto_L1642 := true;
                        end if;
                        goto_L1642 := goto_L1642;
                      end if;
                      goto_L1642 := goto_L1642;
                      if (NOT goto_L1642) then
                        null; -- label L1652
                        -- got s@AO in r1635
                        r1653 := rewire_r1_969(r1635);
                        r1641 := r1653;
                        goto_L1642 := true;
                      end if;
                      goto_L1642 := goto_L1642;
                    end if;
                    goto_L1642 := goto_L1642;
                    if (NOT goto_L1642) then
                      null; -- label L1645
                      -- got s@AO in r1635
                      r1646 := rewire_r0_930(r1635);
                      r1641 := r1646;
                      goto_L1642 := true;
                    end if;
                    goto_L1642 := goto_L1642;
                    null; -- label L1642
                    -- end case
                    r1669 := statevar0;
                    -- got s@AQ in r1669
                    r1672 := rewire_outputs_144(r1669);
                    r1674 := statevar0;
                    -- got s@AS in r1674
                    -- got o@AR in r1672
                    r1678 := "1";
                    r1680 := rewire_setWeOut_853(r1672,r1678);
                    r1682 := rewire_setOutputs_91(r1674,r1680);
                    statevar0 := r1682;
                    r1685 := statevar0;
                    -- got s@AU in r1685
                    r1688 := rewire_outputs_144(r1685);
                    r1690 := statevar0;
                    -- got s@B0 in r1690
                    -- got o@AV in r1688
                    -- got v@AP in r1641
                    r1695 := rewire_setDataOut_1090(r1688,r1641);
                    r1697 := rewire_setOutputs_91(r1690,r1695);
                    statevar0 := r1697;
                    r1700 := statevar0;
                    -- got s@B2 in r1700
                    r1703 := rewire_outputs_144(r1700);
                    r1705 := statevar0;
                    -- got s@B4 in r1705
                    -- got o@B3 in r1703
                    -- got a@AN in r1607
                    r1710 := rewire_setAddrOut_782(r1703,r1607);
                    r1712 := rewire_setOutputs_91(r1705,r1710);
                    statevar0 := r1712;
                    r1715 := statevar0;
                    -- got s@B6 in r1715
                    r1718 := rewire_outputs_144(r1715);
                    -- got o@B7 in r1718
                    nextout := r1718;
                    state := STATE1723;
                    goto_L5439 := true;
                  end if;
                  goto_L5439 := goto_L5439;
                end if;
                goto_L5439 := goto_L5439;
                if (NOT goto_L5439) then
                  null; -- label L1434
                  r1433 := statevar0;
                  -- got c0@9T in r1411
                  -- got c1@9U in r1413
                  r1437 := rewire_mkReg_883(r1411,r1413);
                  b1441 := ("00" = r1437(0 to 1));
                  goto_L1443 := b1441;
                  if (NOT goto_L1443) then
                    goto_L1447 := (NOT b1441);
                    null; -- label L1447
                    -- alt exit (no match)
                    b1448 := ("01" = r1437(0 to 1));
                    goto_L1450 := b1448;
                    if (NOT goto_L1450) then
                      goto_L1454 := (NOT b1448);
                      null; -- label L1454
                      -- alt exit (no match)
                      b1455 := ("10" = r1437(0 to 1));
                      goto_L1457 := b1455;
                      if (NOT goto_L1457) then
                        goto_L1461 := (NOT b1455);
                        null; -- label L1461
                        -- alt exit (no match)
                        -- final pat
                        -- got s@9V in r1433
                        r1464 := rewire_r3_1046(r1433);
                        r1439 := r1464;
                        goto_L1440 := true;
                      end if;
                      goto_L1440 := goto_L1440;
                      if (NOT goto_L1440) then
                        null; -- label L1457
                        -- got s@9V in r1433
                        r1458 := rewire_r2_1008(r1433);
                        r1439 := r1458;
                        goto_L1440 := true;
                      end if;
                      goto_L1440 := goto_L1440;
                    end if;
                    goto_L1440 := goto_L1440;
                    if (NOT goto_L1440) then
                      null; -- label L1450
                      -- got s@9V in r1433
                      r1451 := rewire_r1_969(r1433);
                      r1439 := r1451;
                      goto_L1440 := true;
                    end if;
                    goto_L1440 := goto_L1440;
                  end if;
                  goto_L1440 := goto_L1440;
                  if (NOT goto_L1440) then
                    null; -- label L1443
                    -- got s@9V in r1433
                    r1444 := rewire_r0_930(r1433);
                    r1439 := r1444;
                    goto_L1440 := true;
                  end if;
                  goto_L1440 := goto_L1440;
                  null; -- label L1440
                  -- end case
                  r1467 := statevar0;
                  -- got s@A1 in r1467
                  r1470 := rewire_outputs_144(r1467);
                  r1472 := statevar0;
                  -- got s@A3 in r1472
                  -- got o@A2 in r1470
                  r1476 := "0";
                  r1478 := rewire_setWeOut_853(r1470,r1476);
                  r1480 := rewire_setOutputs_91(r1472,r1478);
                  statevar0 := r1480;
                  r1483 := statevar0;
                  -- got s@A5 in r1483
                  r1486 := rewire_outputs_144(r1483);
                  r1488 := statevar0;
                  -- got s@A7 in r1488
                  -- got o@A6 in r1486
                  -- got a@A0 in r1439
                  r1493 := rewire_setAddrOut_782(r1486,r1439);
                  r1495 := rewire_setOutputs_91(r1488,r1493);
                  statevar0 := r1495;
                  r1498 := statevar0;
                  -- got s@A9 in r1498
                  r1501 := rewire_outputs_144(r1498);
                  -- got o@AA in r1501
                  nextout := r1501;
                  state := STATE1506;
                  goto_L5439 := true;
                end if;
                goto_L5439 := goto_L5439;
              end if;
              goto_L5439 := goto_L5439;
              if (NOT goto_L5439) then
                null; -- label L770
                r769 := statevar0;
                -- got s@8H in r769
                r772 := rewire_pc_462(r769);
                r774 := statevar0;
                -- got s@8J in r774
                r777 := rewire_outputs_144(r774);
                r779 := statevar0;
                -- got s@8L in r779
                -- got o@8K in r777
                -- got pc@8I in r772
                r801 := rewire_setAddrOut_782(r777,r772);
                r803 := rewire_setOutputs_91(r779,r801);
                statevar0 := r803;
                r806 := statevar0;
                -- got s@8N in r806
                r809 := rewire_outputs_144(r806);
                -- got o@8O in r809
                nextout := r809;
                state := STATE814;
                goto_L5439 := true;
              end if;
              goto_L5439 := goto_L5439;
            end if;
            goto_L5439 := goto_L5439;
            if (NOT goto_L5439) then
              null; -- label L418
              r417 := statevar0;
              -- got s@7R in r417
              r455 := "0";
              r457 := rewire_setIEFlag_419(r417,r455);
              statevar0 := r457;
              r460 := statevar0;
              -- got s@7T in r460
              r495 := rewire_pc_462(r460);
              r497 := statevar0;
              -- got s@7V in r497
              r532 := rewire_zFlag_499(r497);
              r534 := statevar0;
              -- got s@81 in r534
              r569 := rewire_cFlag_536(r534);
              r571 := statevar0;
              -- got s@83 in r571
              -- got pc@7U in r495
              r610 := rewire_setPCSave_573(r571,r495);
              statevar0 := r610;
              r613 := statevar0;
              -- got s@85 in r613
              -- got z@80 in r532
              r652 := rewire_setZSave_615(r613,r532);
              statevar0 := r652;
              r655 := statevar0;
              -- got s@87 in r655
              -- got c@82 in r569
              r694 := rewire_setCSave_657(r655,r569);
              statevar0 := r694;
              r697 := statevar0;
              -- got s@89 in r697
              r700 := rewire_outputs_144(r697);
              -- got o@8A in r700
              nextout := r700;
              state := STATE705;
              goto_L5439 := true;
            end if;
            goto_L5439 := goto_L5439;
          end if;
          goto_L5439 := goto_L5439;
          if (NOT goto_L5439) then
            null; -- label L283
            r282 := statevar0;
            -- got s@7E in r282
            r285 := "0";
            r287 := rewire_setCFlag_5(r282,r285);
            statevar0 := r287;
            r290 := statevar0;
            -- got s@7G in r290
            r293 := "0";
            r295 := rewire_setZFlag_48(r290,r293);
            statevar0 := r295;
            r298 := statevar0;
            -- got s@7I in r298
            r301 := rewire_initOutputs_127;
            r303 := rewire_setOutputs_91(r298,r301);
            statevar0 := r303;
            r306 := statevar0;
            -- got s@7K in r306
            r309 := rewire_outputs_144(r306);
            -- got o@7L in r309
            nextout := r309;
            state := STATE314;
            goto_L5439 := true;
          end if;
          goto_L5439 := goto_L5439;
        end if;
        goto_L5439 := goto_L5439;
      end if;
      goto_L5439 := goto_L5439;
      if (NOT goto_L5439) then
        null; -- label L0
        -- START
        -- begin in
        r3 := statevar0;
        -- got s@N2 in r3
        r41 := "0";
        r43 := rewire_setCFlag_5(r3,r41);
        statevar0 := r43;
        r46 := statevar0;
        -- got s@N4 in r46
        r84 := "0";
        r86 := rewire_setZFlag_48(r46,r84);
        statevar0 := r86;
        r89 := statevar0;
        -- got s@N6 in r89
        r137 := rewire_initOutputs_127;
        r139 := rewire_setOutputs_91(r89,r137);
        statevar0 := r139;
        r142 := statevar0;
        -- got s@N8 in r142
        r177 := rewire_outputs_144(r142);
        -- got o@N9 in r177
        nextout := r177;
        state := STATE182;
        goto_L5439 := true;
      end if;
      goto_L5439 := goto_L5439;
      null; -- label L5439
      -- EXIT
    end if;
  end process;
end behavioral;
library ieee;
use ieee.std_logic_1164.all;
-- Uncomment the following line if VHDL primitives are in use.
use work.prims.all;
entity main is
  Port ( clk : in std_logic ;
         input : in std_logic_vector (0 to 9);
         output : out std_logic_vector (0 to 17));
end main;
architecture structural of main is
begin
  dev : entity work.rwcomp0(behavioral)
    port map (clk,input,output);


end structural;
