library ieee;
use ieee.std_logic_1164.all;
-- Uncomment the following line if VHDL primitives are in use.
-- use prims.all;
entity rwcomp0 is
  Port ( clk : in std_logic ;
         input : in std_logic_vector (0 to 895);
         output : out std_logic_vector (0 to 511));
end rwcomp0;

architecture behavioral of rwcomp0 is
  type control_state is (STATE0,STATE1163,STATE2959);
  function rewire_buildSalsa256_1190(r1191 : std_logic_vector ; r1192 : std_logic_vector ; r1193 : std_logic_vector ; r1194 : std_logic_vector) return std_logic_vector;
  function rewire_salsaHash_1666(r1667 : std_logic_vector) return std_logic_vector;
  function rewire_impwords_2610(r2611 : std_logic_vector) return std_logic_vector;
  function rewire_littleendian_2744(r2745 : std_logic_vector) return std_logic_vector;
  function rewire_w8to16le_2839(r2840 : std_logic_vector ; r2841 : std_logic_vector) return std_logic_vector;
  function rewire_w16tow32le_2758(r2759 : std_logic_vector ; r2760 : std_logic_vector) return std_logic_vector;
  function rewire_salsaHashp_1986(r1987 : std_logic_vector) return std_logic_vector;
  function rewire_doubleRound_2024(r2025 : std_logic_vector) return std_logic_vector;
  function rewire_columnRound_2444(r2445 : std_logic_vector) return std_logic_vector;
  function rewire_rowRound_2027(r2028 : std_logic_vector) return std_logic_vector;
  function rewire_quarterRound_2065(r2066 : std_logic_vector) return std_logic_vector;
  function rewire_rot18_2304(r2305 : std_logic_vector) return std_logic_vector;
  function rewire_rot13_2229(r2230 : std_logic_vector) return std_logic_vector;
  function rewire_rot9_2154(r2155 : std_logic_vector) return std_logic_vector;
  function rewire_rot7_2079(r2080 : std_logic_vector) return std_logic_vector;
  function rewire_expwords_1669(r1670 : std_logic_vector) return std_logic_vector;
  function rewire_littleendianp_1707(r1708 : std_logic_vector) return std_logic_vector;
  function rewire_sigma3_1541 return std_logic_vector;
  function rewire_sigma2_1464 return std_logic_vector;
  function rewire_sigma1_1387 return std_logic_vector;
  function rewire_sigma0_1310 return std_logic_vector;
  function rewire_zerothoutput_3 return std_logic_vector;

  function rewire_buildSalsa256_1190(r1191 : std_logic_vector ; r1192 : std_logic_vector ; r1193 : std_logic_vector ; r1194 : std_logic_vector) return std_logic_vector
  is
    variable r2946 : std_logic_vector(0 to 511) := (others => '0');
    variable r2945 : std_logic_vector(0 to 511) := (others => '0');
    variable r1668 : std_logic_vector(0 to 511) := (others => '0');
    variable r1667 : std_logic_vector(0 to 511) := (others => '0');
    variable b1665 : boolean := false;
    variable b1664 : boolean := false;
    variable b1663 : boolean := false;
    variable b1662 : boolean := false;
    variable b1661 : boolean := false;
    variable b1660 : boolean := false;
    variable r1659 : std_logic_vector(0 to 7) := (others => '0');
    variable r1658 : std_logic_vector(0 to 7) := (others => '0');
    variable r1657 : std_logic_vector(0 to 7) := (others => '0');
    variable r1656 : std_logic_vector(0 to 7) := (others => '0');
    variable b1655 : boolean := false;
    variable b1654 : boolean := false;
    variable b1653 : boolean := false;
    variable b1652 : boolean := false;
    variable b1651 : boolean := false;
    variable b1650 : boolean := false;
    variable r1649 : std_logic_vector(0 to 7) := (others => '0');
    variable r1648 : std_logic_vector(0 to 7) := (others => '0');
    variable r1647 : std_logic_vector(0 to 7) := (others => '0');
    variable r1646 : std_logic_vector(0 to 7) := (others => '0');
    variable b1645 : boolean := false;
    variable b1644 : boolean := false;
    variable b1643 : boolean := false;
    variable b1642 : boolean := false;
    variable b1641 : boolean := false;
    variable b1640 : boolean := false;
    variable r1639 : std_logic_vector(0 to 7) := (others => '0');
    variable r1638 : std_logic_vector(0 to 7) := (others => '0');
    variable r1637 : std_logic_vector(0 to 7) := (others => '0');
    variable r1636 : std_logic_vector(0 to 7) := (others => '0');
    variable b1635 : boolean := false;
    variable b1634 : boolean := false;
    variable b1633 : boolean := false;
    variable b1632 : boolean := false;
    variable b1631 : boolean := false;
    variable b1630 : boolean := false;
    variable r1629 : std_logic_vector(0 to 7) := (others => '0');
    variable r1628 : std_logic_vector(0 to 7) := (others => '0');
    variable r1627 : std_logic_vector(0 to 7) := (others => '0');
    variable r1626 : std_logic_vector(0 to 7) := (others => '0');
    variable b1625 : boolean := false;
    variable r1624 : std_logic_vector(0 to 31) := (others => '0');
    variable r1623 : std_logic_vector(0 to 31) := (others => '0');
    variable r1622 : std_logic_vector(0 to 31) := (others => '0');
    variable r1621 : std_logic_vector(0 to 31) := (others => '0');
    variable b1620 : boolean := false;
    variable r1619 : std_logic_vector(0 to 511) := (others => '0');
    variable r1618 : std_logic_vector(0 to 127) := (others => '0');
    variable r1617 : std_logic_vector(0 to 31) := (others => '0');
    variable r1542 : std_logic_vector(0 to 31) := (others => '0');
    variable r1540 : std_logic_vector(0 to 31) := (others => '0');
    variable r1465 : std_logic_vector(0 to 31) := (others => '0');
    variable r1463 : std_logic_vector(0 to 31) := (others => '0');
    variable r1388 : std_logic_vector(0 to 31) := (others => '0');
    variable r1386 : std_logic_vector(0 to 31) := (others => '0');
    variable r1311 : std_logic_vector(0 to 31) := (others => '0');
    variable b1308 : boolean := false;
    variable b1307 : boolean := false;
    variable b1306 : boolean := false;
    variable b1305 : boolean := false;
    variable b1304 : boolean := false;
    variable b1303 : boolean := false;
    variable b1302 : boolean := false;
    variable b1301 : boolean := false;
    variable b1300 : boolean := false;
    variable b1299 : boolean := false;
    variable r1298 : std_logic_vector(0 to 7) := (others => '0');
    variable r1297 : std_logic_vector(0 to 7) := (others => '0');
    variable r1296 : std_logic_vector(0 to 7) := (others => '0');
    variable r1295 : std_logic_vector(0 to 7) := (others => '0');
    variable r1294 : std_logic_vector(0 to 7) := (others => '0');
    variable r1293 : std_logic_vector(0 to 7) := (others => '0');
    variable r1292 : std_logic_vector(0 to 7) := (others => '0');
    variable r1291 : std_logic_vector(0 to 7) := (others => '0');
    variable b1290 : boolean := false;
    variable b1289 : boolean := false;
    variable b1288 : boolean := false;
    variable b1287 : boolean := false;
    variable b1286 : boolean := false;
    variable b1285 : boolean := false;
    variable b1284 : boolean := false;
    variable b1283 : boolean := false;
    variable b1282 : boolean := false;
    variable b1281 : boolean := false;
    variable r1280 : std_logic_vector(0 to 7) := (others => '0');
    variable r1279 : std_logic_vector(0 to 7) := (others => '0');
    variable r1278 : std_logic_vector(0 to 7) := (others => '0');
    variable r1277 : std_logic_vector(0 to 7) := (others => '0');
    variable r1276 : std_logic_vector(0 to 7) := (others => '0');
    variable r1275 : std_logic_vector(0 to 7) := (others => '0');
    variable r1274 : std_logic_vector(0 to 7) := (others => '0');
    variable r1273 : std_logic_vector(0 to 7) := (others => '0');
    variable b1272 : boolean := false;
    variable b1271 : boolean := false;
    variable b1270 : boolean := false;
    variable b1269 : boolean := false;
    variable b1268 : boolean := false;
    variable b1267 : boolean := false;
    variable b1266 : boolean := false;
    variable b1265 : boolean := false;
    variable b1264 : boolean := false;
    variable b1263 : boolean := false;
    variable b1262 : boolean := false;
    variable b1261 : boolean := false;
    variable b1260 : boolean := false;
    variable b1259 : boolean := false;
    variable b1258 : boolean := false;
    variable b1257 : boolean := false;
    variable b1256 : boolean := false;
    variable b1255 : boolean := false;
    variable r1254 : std_logic_vector(0 to 7) := (others => '0');
    variable r1253 : std_logic_vector(0 to 7) := (others => '0');
    variable r1252 : std_logic_vector(0 to 7) := (others => '0');
    variable r1251 : std_logic_vector(0 to 7) := (others => '0');
    variable r1250 : std_logic_vector(0 to 7) := (others => '0');
    variable r1249 : std_logic_vector(0 to 7) := (others => '0');
    variable r1248 : std_logic_vector(0 to 7) := (others => '0');
    variable r1247 : std_logic_vector(0 to 7) := (others => '0');
    variable r1246 : std_logic_vector(0 to 7) := (others => '0');
    variable r1245 : std_logic_vector(0 to 7) := (others => '0');
    variable r1244 : std_logic_vector(0 to 7) := (others => '0');
    variable r1243 : std_logic_vector(0 to 7) := (others => '0');
    variable r1242 : std_logic_vector(0 to 7) := (others => '0');
    variable r1241 : std_logic_vector(0 to 7) := (others => '0');
    variable r1240 : std_logic_vector(0 to 7) := (others => '0');
    variable r1239 : std_logic_vector(0 to 7) := (others => '0');
    variable b1238 : boolean := false;
    variable b1237 : boolean := false;
    variable b1236 : boolean := false;
    variable b1235 : boolean := false;
    variable b1234 : boolean := false;
    variable b1233 : boolean := false;
    variable b1232 : boolean := false;
    variable b1231 : boolean := false;
    variable b1230 : boolean := false;
    variable b1229 : boolean := false;
    variable b1228 : boolean := false;
    variable b1227 : boolean := false;
    variable b1226 : boolean := false;
    variable b1225 : boolean := false;
    variable b1224 : boolean := false;
    variable b1223 : boolean := false;
    variable b1222 : boolean := false;
    variable b1221 : boolean := false;
    variable r1220 : std_logic_vector(0 to 7) := (others => '0');
    variable r1219 : std_logic_vector(0 to 7) := (others => '0');
    variable r1218 : std_logic_vector(0 to 7) := (others => '0');
    variable r1217 : std_logic_vector(0 to 7) := (others => '0');
    variable r1216 : std_logic_vector(0 to 7) := (others => '0');
    variable r1215 : std_logic_vector(0 to 7) := (others => '0');
    variable r1214 : std_logic_vector(0 to 7) := (others => '0');
    variable r1213 : std_logic_vector(0 to 7) := (others => '0');
    variable r1212 : std_logic_vector(0 to 7) := (others => '0');
    variable r1211 : std_logic_vector(0 to 7) := (others => '0');
    variable r1210 : std_logic_vector(0 to 7) := (others => '0');
    variable r1209 : std_logic_vector(0 to 7) := (others => '0');
    variable r1208 : std_logic_vector(0 to 7) := (others => '0');
    variable r1207 : std_logic_vector(0 to 7) := (others => '0');
    variable r1206 : std_logic_vector(0 to 7) := (others => '0');
    variable r1205 : std_logic_vector(0 to 7) := (others => '0');
    variable b1204 : boolean := false;
    variable r1203 : std_logic_vector(0 to 63) := (others => '0');
    variable r1202 : std_logic_vector(0 to 63) := (others => '0');
    variable r1201 : std_logic_vector(0 to 127) := (others => '0');
    variable r1200 : std_logic_vector(0 to 127) := (others => '0');
    variable b1199 : boolean := false;
    variable r1198 : std_logic_vector(0 to 511) := (others => '0');
    variable r1197 : std_logic_vector(0 to 383) := (others => '0');
  begin
    b1199 := true;
    r1200 := r1197(0 to 127);
    r1201 := r1197(128 to 255);
    r1202 := r1197(256 to 319);
    r1203 := r1197(320 to 383);
    b1204 := true;
    r1205 := r1200(0 to 7);
    r1206 := r1200(8 to 15);
    r1207 := r1200(16 to 23);
    r1208 := r1200(24 to 31);
    r1209 := r1200(32 to 39);
    r1210 := r1200(40 to 47);
    r1211 := r1200(48 to 55);
    r1212 := r1200(56 to 63);
    r1213 := r1200(64 to 71);
    r1214 := r1200(72 to 79);
    r1215 := r1200(80 to 87);
    r1216 := r1200(88 to 95);
    r1217 := r1200(96 to 103);
    r1218 := r1200(104 to 111);
    r1219 := r1200(112 to 119);
    r1220 := r1200(120 to 127);
    b1221 := true;
    b1222 := true;
    b1223 := true;
    b1224 := true;
    b1225 := true;
    b1226 := true;
    b1227 := true;
    b1228 := true;
    b1229 := true;
    b1230 := true;
    b1231 := true;
    b1232 := true;
    b1233 := true;
    b1234 := true;
    b1235 := true;
    b1236 := true;
    b1237 := (b1221 AND (b1222 AND (b1223 AND (b1224 AND (b1225 AND (b1226 AND (b1227 AND (b1228 AND (b1229 AND (b1230 AND (b1231 AND (b1232 AND (b1233 AND (b1234 AND (b1235 AND b1236)))))))))))))));
    b1238 := true;
    r1239 := r1201(0 to 7);
    r1240 := r1201(8 to 15);
    r1241 := r1201(16 to 23);
    r1242 := r1201(24 to 31);
    r1243 := r1201(32 to 39);
    r1244 := r1201(40 to 47);
    r1245 := r1201(48 to 55);
    r1246 := r1201(56 to 63);
    r1247 := r1201(64 to 71);
    r1248 := r1201(72 to 79);
    r1249 := r1201(80 to 87);
    r1250 := r1201(88 to 95);
    r1251 := r1201(96 to 103);
    r1252 := r1201(104 to 111);
    r1253 := r1201(112 to 119);
    r1254 := r1201(120 to 127);
    b1255 := true;
    b1256 := true;
    b1257 := true;
    b1258 := true;
    b1259 := true;
    b1260 := true;
    b1261 := true;
    b1262 := true;
    b1263 := true;
    b1264 := true;
    b1265 := true;
    b1266 := true;
    b1267 := true;
    b1268 := true;
    b1269 := true;
    b1270 := true;
    b1271 := (b1255 AND (b1256 AND (b1257 AND (b1258 AND (b1259 AND (b1260 AND (b1261 AND (b1262 AND (b1263 AND (b1264 AND (b1265 AND (b1266 AND (b1267 AND (b1268 AND (b1269 AND b1270)))))))))))))));
    b1272 := true;
    r1273 := r1202(0 to 7);
    r1274 := r1202(8 to 15);
    r1275 := r1202(16 to 23);
    r1276 := r1202(24 to 31);
    r1277 := r1202(32 to 39);
    r1278 := r1202(40 to 47);
    r1279 := r1202(48 to 55);
    r1280 := r1202(56 to 63);
    b1281 := true;
    b1282 := true;
    b1283 := true;
    b1284 := true;
    b1285 := true;
    b1286 := true;
    b1287 := true;
    b1288 := true;
    b1289 := (b1281 AND (b1282 AND (b1283 AND (b1284 AND (b1285 AND (b1286 AND (b1287 AND b1288)))))));
    b1290 := true;
    r1291 := r1203(0 to 7);
    r1292 := r1203(8 to 15);
    r1293 := r1203(16 to 23);
    r1294 := r1203(24 to 31);
    r1295 := r1203(32 to 39);
    r1296 := r1203(40 to 47);
    r1297 := r1203(48 to 55);
    r1298 := r1203(56 to 63);
    b1299 := true;
    b1300 := true;
    b1301 := true;
    b1302 := true;
    b1303 := true;
    b1304 := true;
    b1305 := true;
    b1306 := true;
    b1307 := (b1299 AND (b1300 AND (b1301 AND (b1302 AND (b1303 AND (b1304 AND (b1305 AND b1306)))))));
    b1308 := (b1237 AND (b1271 AND (b1289 AND b1307)));
    if b1308 then
      b1620 := true;
      r1621 := r1618(0 to 31);
      r1622 := r1618(32 to 63);
      r1623 := r1618(64 to 95);
      r1624 := r1618(96 to 127);
      b1625 := true;
      r1626 := r1621(0 to 7);
      r1627 := r1621(8 to 15);
      r1628 := r1621(16 to 23);
      r1629 := r1621(24 to 31);
      b1630 := true;
      b1631 := true;
      b1632 := true;
      b1633 := true;
      b1634 := (b1630 AND (b1631 AND (b1632 AND b1633)));
      b1635 := true;
      r1636 := r1622(0 to 7);
      r1637 := r1622(8 to 15);
      r1638 := r1622(16 to 23);
      r1639 := r1622(24 to 31);
      b1640 := true;
      b1641 := true;
      b1642 := true;
      b1643 := true;
      b1644 := (b1640 AND (b1641 AND (b1642 AND b1643)));
      b1645 := true;
      r1646 := r1623(0 to 7);
      r1647 := r1623(8 to 15);
      r1648 := r1623(16 to 23);
      r1649 := r1623(24 to 31);
      b1650 := true;
      b1651 := true;
      b1652 := true;
      b1653 := true;
      b1654 := (b1650 AND (b1651 AND (b1652 AND b1653)));
      b1655 := true;
      r1656 := r1624(0 to 7);
      r1657 := r1624(8 to 15);
      r1658 := r1624(16 to 23);
      r1659 := r1624(24 to 31);
      b1660 := true;
      b1661 := true;
      b1662 := true;
      b1663 := true;
      b1664 := (b1660 AND (b1661 AND (b1662 AND b1663)));
      b1665 := (b1634 AND (b1644 AND (b1654 AND b1664)));
      if b1665 then
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        r2945 := (r1626 & r1627 & r1628 & r1629 & r1205 & r1206 & r1207 & r1208 & r1209 & r1210 & r1211 & r1212 & r1213 & r1214 & r1215 & r1216 & r1217 & r1218 & r1219 & r1220 & r1636 & r1637 & r1638 & r1639 & r1273 & r1274 & r1275 & r1276 & r1277 & r1278 & r1279 & r1280 & r1291 & r1292 & r1293 & r1294 & r1295 & r1296 & r1297 & r1298 & r1646 & r1647 & r1648 & r1649 & r1239 & r1240 & r1241 & r1242 & r1243 & r1244 & r1245 & r1246 & r1247 & r1248 & r1249 & r1250 & r1251 & r1252 & r1253 & r1254 & r1656 & r1657 & r1658 & r1659);
        r2946 := rewire_salsaHash_1666(r2945);
        r1619 := r2946;
      end if;
      r1198 := r1619;
    end if;
    return r1198;
  end rewire_buildSalsa256_1190;
  function rewire_salsaHash_1666(r1667 : std_logic_vector) return std_logic_vector
  is
    variable r2943 : std_logic_vector(0 to 511) := (others => '0');
    variable r2942 : std_logic_vector(0 to 511) := (others => '0');
    variable r2941 : std_logic_vector(0 to 511) := (others => '0');
    variable r2612 : std_logic_vector(0 to 511) := (others => '0');
    variable r2611 : std_logic_vector(0 to 511) := (others => '0');
    variable r1988 : std_logic_vector(0 to 511) := (others => '0');
    variable r1987 : std_logic_vector(0 to 511) := (others => '0');
    variable r1671 : std_logic_vector(0 to 511) := (others => '0');
    variable r1670 : std_logic_vector(0 to 511) := (others => '0');
  begin
    null;
    r2941 := rewire_impwords_2610(r1667);
    r2942 := rewire_salsaHashp_1986(r2941);
    r2943 := rewire_expwords_1669(r2942);
    return r2943;
  end rewire_salsaHash_1666;
  function rewire_impwords_2610(r2611 : std_logic_vector) return std_logic_vector
  is
    variable r2940 : std_logic_vector(0 to 511) := (others => '0');
    variable r2938 : std_logic_vector(0 to 31) := (others => '0');
    variable r2937 : std_logic_vector(0 to 31) := (others => '0');
    variable r2935 : std_logic_vector(0 to 31) := (others => '0');
    variable r2934 : std_logic_vector(0 to 31) := (others => '0');
    variable r2932 : std_logic_vector(0 to 31) := (others => '0');
    variable r2931 : std_logic_vector(0 to 31) := (others => '0');
    variable r2929 : std_logic_vector(0 to 31) := (others => '0');
    variable r2928 : std_logic_vector(0 to 31) := (others => '0');
    variable r2926 : std_logic_vector(0 to 31) := (others => '0');
    variable r2925 : std_logic_vector(0 to 31) := (others => '0');
    variable r2923 : std_logic_vector(0 to 31) := (others => '0');
    variable r2922 : std_logic_vector(0 to 31) := (others => '0');
    variable r2920 : std_logic_vector(0 to 31) := (others => '0');
    variable r2919 : std_logic_vector(0 to 31) := (others => '0');
    variable r2917 : std_logic_vector(0 to 31) := (others => '0');
    variable r2916 : std_logic_vector(0 to 31) := (others => '0');
    variable r2914 : std_logic_vector(0 to 31) := (others => '0');
    variable r2913 : std_logic_vector(0 to 31) := (others => '0');
    variable r2911 : std_logic_vector(0 to 31) := (others => '0');
    variable r2910 : std_logic_vector(0 to 31) := (others => '0');
    variable r2908 : std_logic_vector(0 to 31) := (others => '0');
    variable r2907 : std_logic_vector(0 to 31) := (others => '0');
    variable r2905 : std_logic_vector(0 to 31) := (others => '0');
    variable r2904 : std_logic_vector(0 to 31) := (others => '0');
    variable r2902 : std_logic_vector(0 to 31) := (others => '0');
    variable r2901 : std_logic_vector(0 to 31) := (others => '0');
    variable r2899 : std_logic_vector(0 to 31) := (others => '0');
    variable r2898 : std_logic_vector(0 to 31) := (others => '0');
    variable r2896 : std_logic_vector(0 to 31) := (others => '0');
    variable r2895 : std_logic_vector(0 to 31) := (others => '0');
    variable r2893 : std_logic_vector(0 to 31) := (others => '0');
    variable r2892 : std_logic_vector(0 to 31) := (others => '0');
    variable r2746 : std_logic_vector(0 to 31) := (others => '0');
    variable r2745 : std_logic_vector(0 to 31) := (others => '0');
    variable b2743 : boolean := false;
    variable b2742 : boolean := false;
    variable b2741 : boolean := false;
    variable b2740 : boolean := false;
    variable b2739 : boolean := false;
    variable b2738 : boolean := false;
    variable b2737 : boolean := false;
    variable b2736 : boolean := false;
    variable b2735 : boolean := false;
    variable b2734 : boolean := false;
    variable b2733 : boolean := false;
    variable b2732 : boolean := false;
    variable b2731 : boolean := false;
    variable b2730 : boolean := false;
    variable b2729 : boolean := false;
    variable b2728 : boolean := false;
    variable b2727 : boolean := false;
    variable b2726 : boolean := false;
    variable b2725 : boolean := false;
    variable b2724 : boolean := false;
    variable b2723 : boolean := false;
    variable b2722 : boolean := false;
    variable b2721 : boolean := false;
    variable b2720 : boolean := false;
    variable b2719 : boolean := false;
    variable b2718 : boolean := false;
    variable b2717 : boolean := false;
    variable b2716 : boolean := false;
    variable b2715 : boolean := false;
    variable b2714 : boolean := false;
    variable b2713 : boolean := false;
    variable b2712 : boolean := false;
    variable b2711 : boolean := false;
    variable b2710 : boolean := false;
    variable b2709 : boolean := false;
    variable b2708 : boolean := false;
    variable b2707 : boolean := false;
    variable b2706 : boolean := false;
    variable b2705 : boolean := false;
    variable b2704 : boolean := false;
    variable b2703 : boolean := false;
    variable b2702 : boolean := false;
    variable b2701 : boolean := false;
    variable b2700 : boolean := false;
    variable b2699 : boolean := false;
    variable b2698 : boolean := false;
    variable b2697 : boolean := false;
    variable b2696 : boolean := false;
    variable b2695 : boolean := false;
    variable b2694 : boolean := false;
    variable b2693 : boolean := false;
    variable b2692 : boolean := false;
    variable b2691 : boolean := false;
    variable b2690 : boolean := false;
    variable b2689 : boolean := false;
    variable b2688 : boolean := false;
    variable b2687 : boolean := false;
    variable b2686 : boolean := false;
    variable b2685 : boolean := false;
    variable b2684 : boolean := false;
    variable b2683 : boolean := false;
    variable b2682 : boolean := false;
    variable b2681 : boolean := false;
    variable b2680 : boolean := false;
    variable b2679 : boolean := false;
    variable r2678 : std_logic_vector(0 to 7) := (others => '0');
    variable r2677 : std_logic_vector(0 to 7) := (others => '0');
    variable r2676 : std_logic_vector(0 to 7) := (others => '0');
    variable r2675 : std_logic_vector(0 to 7) := (others => '0');
    variable r2674 : std_logic_vector(0 to 7) := (others => '0');
    variable r2673 : std_logic_vector(0 to 7) := (others => '0');
    variable r2672 : std_logic_vector(0 to 7) := (others => '0');
    variable r2671 : std_logic_vector(0 to 7) := (others => '0');
    variable r2670 : std_logic_vector(0 to 7) := (others => '0');
    variable r2669 : std_logic_vector(0 to 7) := (others => '0');
    variable r2668 : std_logic_vector(0 to 7) := (others => '0');
    variable r2667 : std_logic_vector(0 to 7) := (others => '0');
    variable r2666 : std_logic_vector(0 to 7) := (others => '0');
    variable r2665 : std_logic_vector(0 to 7) := (others => '0');
    variable r2664 : std_logic_vector(0 to 7) := (others => '0');
    variable r2663 : std_logic_vector(0 to 7) := (others => '0');
    variable r2662 : std_logic_vector(0 to 7) := (others => '0');
    variable r2661 : std_logic_vector(0 to 7) := (others => '0');
    variable r2660 : std_logic_vector(0 to 7) := (others => '0');
    variable r2659 : std_logic_vector(0 to 7) := (others => '0');
    variable r2658 : std_logic_vector(0 to 7) := (others => '0');
    variable r2657 : std_logic_vector(0 to 7) := (others => '0');
    variable r2656 : std_logic_vector(0 to 7) := (others => '0');
    variable r2655 : std_logic_vector(0 to 7) := (others => '0');
    variable r2654 : std_logic_vector(0 to 7) := (others => '0');
    variable r2653 : std_logic_vector(0 to 7) := (others => '0');
    variable r2652 : std_logic_vector(0 to 7) := (others => '0');
    variable r2651 : std_logic_vector(0 to 7) := (others => '0');
    variable r2650 : std_logic_vector(0 to 7) := (others => '0');
    variable r2649 : std_logic_vector(0 to 7) := (others => '0');
    variable r2648 : std_logic_vector(0 to 7) := (others => '0');
    variable r2647 : std_logic_vector(0 to 7) := (others => '0');
    variable r2646 : std_logic_vector(0 to 7) := (others => '0');
    variable r2645 : std_logic_vector(0 to 7) := (others => '0');
    variable r2644 : std_logic_vector(0 to 7) := (others => '0');
    variable r2643 : std_logic_vector(0 to 7) := (others => '0');
    variable r2642 : std_logic_vector(0 to 7) := (others => '0');
    variable r2641 : std_logic_vector(0 to 7) := (others => '0');
    variable r2640 : std_logic_vector(0 to 7) := (others => '0');
    variable r2639 : std_logic_vector(0 to 7) := (others => '0');
    variable r2638 : std_logic_vector(0 to 7) := (others => '0');
    variable r2637 : std_logic_vector(0 to 7) := (others => '0');
    variable r2636 : std_logic_vector(0 to 7) := (others => '0');
    variable r2635 : std_logic_vector(0 to 7) := (others => '0');
    variable r2634 : std_logic_vector(0 to 7) := (others => '0');
    variable r2633 : std_logic_vector(0 to 7) := (others => '0');
    variable r2632 : std_logic_vector(0 to 7) := (others => '0');
    variable r2631 : std_logic_vector(0 to 7) := (others => '0');
    variable r2630 : std_logic_vector(0 to 7) := (others => '0');
    variable r2629 : std_logic_vector(0 to 7) := (others => '0');
    variable r2628 : std_logic_vector(0 to 7) := (others => '0');
    variable r2627 : std_logic_vector(0 to 7) := (others => '0');
    variable r2626 : std_logic_vector(0 to 7) := (others => '0');
    variable r2625 : std_logic_vector(0 to 7) := (others => '0');
    variable r2624 : std_logic_vector(0 to 7) := (others => '0');
    variable r2623 : std_logic_vector(0 to 7) := (others => '0');
    variable r2622 : std_logic_vector(0 to 7) := (others => '0');
    variable r2621 : std_logic_vector(0 to 7) := (others => '0');
    variable r2620 : std_logic_vector(0 to 7) := (others => '0');
    variable r2619 : std_logic_vector(0 to 7) := (others => '0');
    variable r2618 : std_logic_vector(0 to 7) := (others => '0');
    variable r2617 : std_logic_vector(0 to 7) := (others => '0');
    variable r2616 : std_logic_vector(0 to 7) := (others => '0');
    variable r2615 : std_logic_vector(0 to 7) := (others => '0');
    variable b2614 : boolean := false;
    variable r2613 : std_logic_vector(0 to 511) := (others => '0');
  begin
    b2614 := true;
    r2615 := r2611(0 to 7);
    r2616 := r2611(8 to 15);
    r2617 := r2611(16 to 23);
    r2618 := r2611(24 to 31);
    r2619 := r2611(32 to 39);
    r2620 := r2611(40 to 47);
    r2621 := r2611(48 to 55);
    r2622 := r2611(56 to 63);
    r2623 := r2611(64 to 71);
    r2624 := r2611(72 to 79);
    r2625 := r2611(80 to 87);
    r2626 := r2611(88 to 95);
    r2627 := r2611(96 to 103);
    r2628 := r2611(104 to 111);
    r2629 := r2611(112 to 119);
    r2630 := r2611(120 to 127);
    r2631 := r2611(128 to 135);
    r2632 := r2611(136 to 143);
    r2633 := r2611(144 to 151);
    r2634 := r2611(152 to 159);
    r2635 := r2611(160 to 167);
    r2636 := r2611(168 to 175);
    r2637 := r2611(176 to 183);
    r2638 := r2611(184 to 191);
    r2639 := r2611(192 to 199);
    r2640 := r2611(200 to 207);
    r2641 := r2611(208 to 215);
    r2642 := r2611(216 to 223);
    r2643 := r2611(224 to 231);
    r2644 := r2611(232 to 239);
    r2645 := r2611(240 to 247);
    r2646 := r2611(248 to 255);
    r2647 := r2611(256 to 263);
    r2648 := r2611(264 to 271);
    r2649 := r2611(272 to 279);
    r2650 := r2611(280 to 287);
    r2651 := r2611(288 to 295);
    r2652 := r2611(296 to 303);
    r2653 := r2611(304 to 311);
    r2654 := r2611(312 to 319);
    r2655 := r2611(320 to 327);
    r2656 := r2611(328 to 335);
    r2657 := r2611(336 to 343);
    r2658 := r2611(344 to 351);
    r2659 := r2611(352 to 359);
    r2660 := r2611(360 to 367);
    r2661 := r2611(368 to 375);
    r2662 := r2611(376 to 383);
    r2663 := r2611(384 to 391);
    r2664 := r2611(392 to 399);
    r2665 := r2611(400 to 407);
    r2666 := r2611(408 to 415);
    r2667 := r2611(416 to 423);
    r2668 := r2611(424 to 431);
    r2669 := r2611(432 to 439);
    r2670 := r2611(440 to 447);
    r2671 := r2611(448 to 455);
    r2672 := r2611(456 to 463);
    r2673 := r2611(464 to 471);
    r2674 := r2611(472 to 479);
    r2675 := r2611(480 to 487);
    r2676 := r2611(488 to 495);
    r2677 := r2611(496 to 503);
    r2678 := r2611(504 to 511);
    b2679 := true;
    b2680 := true;
    b2681 := true;
    b2682 := true;
    b2683 := true;
    b2684 := true;
    b2685 := true;
    b2686 := true;
    b2687 := true;
    b2688 := true;
    b2689 := true;
    b2690 := true;
    b2691 := true;
    b2692 := true;
    b2693 := true;
    b2694 := true;
    b2695 := true;
    b2696 := true;
    b2697 := true;
    b2698 := true;
    b2699 := true;
    b2700 := true;
    b2701 := true;
    b2702 := true;
    b2703 := true;
    b2704 := true;
    b2705 := true;
    b2706 := true;
    b2707 := true;
    b2708 := true;
    b2709 := true;
    b2710 := true;
    b2711 := true;
    b2712 := true;
    b2713 := true;
    b2714 := true;
    b2715 := true;
    b2716 := true;
    b2717 := true;
    b2718 := true;
    b2719 := true;
    b2720 := true;
    b2721 := true;
    b2722 := true;
    b2723 := true;
    b2724 := true;
    b2725 := true;
    b2726 := true;
    b2727 := true;
    b2728 := true;
    b2729 := true;
    b2730 := true;
    b2731 := true;
    b2732 := true;
    b2733 := true;
    b2734 := true;
    b2735 := true;
    b2736 := true;
    b2737 := true;
    b2738 := true;
    b2739 := true;
    b2740 := true;
    b2741 := true;
    b2742 := true;
    b2743 := (b2679 AND (b2680 AND (b2681 AND (b2682 AND (b2683 AND (b2684 AND (b2685 AND (b2686 AND (b2687 AND (b2688 AND (b2689 AND (b2690 AND (b2691 AND (b2692 AND (b2693 AND (b2694 AND (b2695 AND (b2696 AND (b2697 AND (b2698 AND (b2699 AND (b2700 AND (b2701 AND (b2702 AND (b2703 AND (b2704 AND (b2705 AND (b2706 AND (b2707 AND (b2708 AND (b2709 AND (b2710 AND (b2711 AND (b2712 AND (b2713 AND (b2714 AND (b2715 AND (b2716 AND (b2717 AND (b2718 AND (b2719 AND (b2720 AND (b2721 AND (b2722 AND (b2723 AND (b2724 AND (b2725 AND (b2726 AND (b2727 AND (b2728 AND (b2729 AND (b2730 AND (b2731 AND (b2732 AND (b2733 AND (b2734 AND (b2735 AND (b2736 AND (b2737 AND (b2738 AND (b2739 AND (b2740 AND (b2741 AND b2742)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
    if b2743 then
      null;
      null;
      null;
      null;
      r2892 := (r2615 & r2616 & r2617 & r2618);
      r2893 := rewire_littleendian_2744(r2892);
      null;
      null;
      null;
      null;
      r2895 := (r2619 & r2620 & r2621 & r2622);
      r2896 := rewire_littleendian_2744(r2895);
      null;
      null;
      null;
      null;
      r2898 := (r2623 & r2624 & r2625 & r2626);
      r2899 := rewire_littleendian_2744(r2898);
      null;
      null;
      null;
      null;
      r2901 := (r2627 & r2628 & r2629 & r2630);
      r2902 := rewire_littleendian_2744(r2901);
      null;
      null;
      null;
      null;
      r2904 := (r2631 & r2632 & r2633 & r2634);
      r2905 := rewire_littleendian_2744(r2904);
      null;
      null;
      null;
      null;
      r2907 := (r2635 & r2636 & r2637 & r2638);
      r2908 := rewire_littleendian_2744(r2907);
      null;
      null;
      null;
      null;
      r2910 := (r2639 & r2640 & r2641 & r2642);
      r2911 := rewire_littleendian_2744(r2910);
      null;
      null;
      null;
      null;
      r2913 := (r2643 & r2644 & r2645 & r2646);
      r2914 := rewire_littleendian_2744(r2913);
      null;
      null;
      null;
      null;
      r2916 := (r2647 & r2648 & r2649 & r2650);
      r2917 := rewire_littleendian_2744(r2916);
      null;
      null;
      null;
      null;
      r2919 := (r2651 & r2652 & r2653 & r2654);
      r2920 := rewire_littleendian_2744(r2919);
      null;
      null;
      null;
      null;
      r2922 := (r2655 & r2656 & r2657 & r2658);
      r2923 := rewire_littleendian_2744(r2922);
      null;
      null;
      null;
      null;
      r2925 := (r2659 & r2660 & r2661 & r2662);
      r2926 := rewire_littleendian_2744(r2925);
      null;
      null;
      null;
      null;
      r2928 := (r2663 & r2664 & r2665 & r2666);
      r2929 := rewire_littleendian_2744(r2928);
      null;
      null;
      null;
      null;
      r2931 := (r2667 & r2668 & r2669 & r2670);
      r2932 := rewire_littleendian_2744(r2931);
      null;
      null;
      null;
      null;
      r2934 := (r2671 & r2672 & r2673 & r2674);
      r2935 := rewire_littleendian_2744(r2934);
      null;
      null;
      null;
      null;
      r2937 := (r2675 & r2676 & r2677 & r2678);
      r2938 := rewire_littleendian_2744(r2937);
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      r2940 := (r2893 & r2896 & r2899 & r2902 & r2905 & r2908 & r2911 & r2914 & r2917 & r2920 & r2923 & r2926 & r2929 & r2932 & r2935 & r2938);
      r2613 := r2940;
    end if;
    return r2613;
  end rewire_impwords_2610;
  function rewire_littleendian_2744(r2745 : std_logic_vector) return std_logic_vector
  is
    variable r2890 : std_logic_vector(0 to 31) := (others => '0');
    variable r2889 : std_logic_vector(0 to 15) := (others => '0');
    variable r2888 : std_logic_vector(0 to 15) := (others => '0');
    variable r2842 : std_logic_vector(0 to 15) := (others => '0');
    variable r2841 : std_logic_vector(0 to 7) := (others => '0');
    variable r2840 : std_logic_vector(0 to 7) := (others => '0');
    variable r2761 : std_logic_vector(0 to 31) := (others => '0');
    variable r2760 : std_logic_vector(0 to 15) := (others => '0');
    variable r2759 : std_logic_vector(0 to 15) := (others => '0');
    variable b2757 : boolean := false;
    variable b2756 : boolean := false;
    variable b2755 : boolean := false;
    variable b2754 : boolean := false;
    variable b2753 : boolean := false;
    variable r2752 : std_logic_vector(0 to 7) := (others => '0');
    variable r2751 : std_logic_vector(0 to 7) := (others => '0');
    variable r2750 : std_logic_vector(0 to 7) := (others => '0');
    variable r2749 : std_logic_vector(0 to 7) := (others => '0');
    variable b2748 : boolean := false;
    variable r2747 : std_logic_vector(0 to 31) := (others => '0');
  begin
    b2748 := true;
    r2749 := r2745(0 to 7);
    r2750 := r2745(8 to 15);
    r2751 := r2745(16 to 23);
    r2752 := r2745(24 to 31);
    b2753 := true;
    b2754 := true;
    b2755 := true;
    b2756 := true;
    b2757 := (b2753 AND (b2754 AND (b2755 AND b2756)));
    if b2757 then
      null;
      null;
      r2888 := rewire_w8to16le_2839(r2752,r2751);
      null;
      null;
      r2889 := rewire_w8to16le_2839(r2750,r2749);
      r2890 := rewire_w16tow32le_2758(r2888,r2889);
      r2747 := r2890;
    end if;
    return r2747;
  end rewire_littleendian_2744;
  function rewire_w8to16le_2839(r2840 : std_logic_vector ; r2841 : std_logic_vector) return std_logic_vector
  is
    variable r2887 : std_logic_vector(0 to 15) := (others => '0');
    variable b2885 : boolean := false;
    variable b2884 : boolean := false;
    variable b2883 : boolean := false;
    variable b2882 : boolean := false;
    variable b2881 : boolean := false;
    variable b2880 : boolean := false;
    variable b2879 : boolean := false;
    variable b2878 : boolean := false;
    variable b2877 : boolean := false;
    variable b2876 : boolean := false;
    variable r2875 : std_logic_vector(0 to 0) := (others => '0');
    variable r2874 : std_logic_vector(0 to 0) := (others => '0');
    variable r2873 : std_logic_vector(0 to 0) := (others => '0');
    variable r2872 : std_logic_vector(0 to 0) := (others => '0');
    variable r2871 : std_logic_vector(0 to 0) := (others => '0');
    variable r2870 : std_logic_vector(0 to 0) := (others => '0');
    variable r2869 : std_logic_vector(0 to 0) := (others => '0');
    variable r2868 : std_logic_vector(0 to 0) := (others => '0');
    variable b2867 : boolean := false;
    variable b2866 : boolean := false;
    variable b2865 : boolean := false;
    variable b2864 : boolean := false;
    variable b2863 : boolean := false;
    variable b2862 : boolean := false;
    variable b2861 : boolean := false;
    variable b2860 : boolean := false;
    variable b2859 : boolean := false;
    variable b2858 : boolean := false;
    variable r2857 : std_logic_vector(0 to 0) := (others => '0');
    variable r2856 : std_logic_vector(0 to 0) := (others => '0');
    variable r2855 : std_logic_vector(0 to 0) := (others => '0');
    variable r2854 : std_logic_vector(0 to 0) := (others => '0');
    variable r2853 : std_logic_vector(0 to 0) := (others => '0');
    variable r2852 : std_logic_vector(0 to 0) := (others => '0');
    variable r2851 : std_logic_vector(0 to 0) := (others => '0');
    variable r2850 : std_logic_vector(0 to 0) := (others => '0');
    variable b2849 : boolean := false;
    variable r2848 : std_logic_vector(0 to 7) := (others => '0');
    variable r2847 : std_logic_vector(0 to 7) := (others => '0');
    variable b2846 : boolean := false;
    variable r2845 : std_logic_vector(0 to 15) := (others => '0');
    variable r2844 : std_logic_vector(0 to 15) := (others => '0');
  begin
    b2846 := true;
    r2847 := r2844(0 to 7);
    r2848 := r2844(8 to 15);
    b2849 := true;
    r2850 := r2847(0 to 0);
    r2851 := r2847(1 to 1);
    r2852 := r2847(2 to 2);
    r2853 := r2847(3 to 3);
    r2854 := r2847(4 to 4);
    r2855 := r2847(5 to 5);
    r2856 := r2847(6 to 6);
    r2857 := r2847(7 to 7);
    b2858 := true;
    b2859 := true;
    b2860 := true;
    b2861 := true;
    b2862 := true;
    b2863 := true;
    b2864 := true;
    b2865 := true;
    b2866 := (b2858 AND (b2859 AND (b2860 AND (b2861 AND (b2862 AND (b2863 AND (b2864 AND b2865)))))));
    b2867 := true;
    r2868 := r2848(0 to 0);
    r2869 := r2848(1 to 1);
    r2870 := r2848(2 to 2);
    r2871 := r2848(3 to 3);
    r2872 := r2848(4 to 4);
    r2873 := r2848(5 to 5);
    r2874 := r2848(6 to 6);
    r2875 := r2848(7 to 7);
    b2876 := true;
    b2877 := true;
    b2878 := true;
    b2879 := true;
    b2880 := true;
    b2881 := true;
    b2882 := true;
    b2883 := true;
    b2884 := (b2876 AND (b2877 AND (b2878 AND (b2879 AND (b2880 AND (b2881 AND (b2882 AND b2883)))))));
    b2885 := (b2866 AND b2884);
    if b2885 then
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      r2887 := (r2868 & r2869 & r2870 & r2871 & r2872 & r2873 & r2874 & r2875 & r2850 & r2851 & r2852 & r2853 & r2854 & r2855 & r2856 & r2857);
      r2845 := r2887;
    end if;
    return r2845;
  end rewire_w8to16le_2839;
  function rewire_w16tow32le_2758(r2759 : std_logic_vector ; r2760 : std_logic_vector) return std_logic_vector
  is
    variable r2838 : std_logic_vector(0 to 31) := (others => '0');
    variable b2836 : boolean := false;
    variable b2835 : boolean := false;
    variable b2834 : boolean := false;
    variable b2833 : boolean := false;
    variable b2832 : boolean := false;
    variable b2831 : boolean := false;
    variable b2830 : boolean := false;
    variable b2829 : boolean := false;
    variable b2828 : boolean := false;
    variable b2827 : boolean := false;
    variable b2826 : boolean := false;
    variable b2825 : boolean := false;
    variable b2824 : boolean := false;
    variable b2823 : boolean := false;
    variable b2822 : boolean := false;
    variable b2821 : boolean := false;
    variable b2820 : boolean := false;
    variable b2819 : boolean := false;
    variable r2818 : std_logic_vector(0 to 0) := (others => '0');
    variable r2817 : std_logic_vector(0 to 0) := (others => '0');
    variable r2816 : std_logic_vector(0 to 0) := (others => '0');
    variable r2815 : std_logic_vector(0 to 0) := (others => '0');
    variable r2814 : std_logic_vector(0 to 0) := (others => '0');
    variable r2813 : std_logic_vector(0 to 0) := (others => '0');
    variable r2812 : std_logic_vector(0 to 0) := (others => '0');
    variable r2811 : std_logic_vector(0 to 0) := (others => '0');
    variable r2810 : std_logic_vector(0 to 0) := (others => '0');
    variable r2809 : std_logic_vector(0 to 0) := (others => '0');
    variable r2808 : std_logic_vector(0 to 0) := (others => '0');
    variable r2807 : std_logic_vector(0 to 0) := (others => '0');
    variable r2806 : std_logic_vector(0 to 0) := (others => '0');
    variable r2805 : std_logic_vector(0 to 0) := (others => '0');
    variable r2804 : std_logic_vector(0 to 0) := (others => '0');
    variable r2803 : std_logic_vector(0 to 0) := (others => '0');
    variable b2802 : boolean := false;
    variable b2801 : boolean := false;
    variable b2800 : boolean := false;
    variable b2799 : boolean := false;
    variable b2798 : boolean := false;
    variable b2797 : boolean := false;
    variable b2796 : boolean := false;
    variable b2795 : boolean := false;
    variable b2794 : boolean := false;
    variable b2793 : boolean := false;
    variable b2792 : boolean := false;
    variable b2791 : boolean := false;
    variable b2790 : boolean := false;
    variable b2789 : boolean := false;
    variable b2788 : boolean := false;
    variable b2787 : boolean := false;
    variable b2786 : boolean := false;
    variable b2785 : boolean := false;
    variable r2784 : std_logic_vector(0 to 0) := (others => '0');
    variable r2783 : std_logic_vector(0 to 0) := (others => '0');
    variable r2782 : std_logic_vector(0 to 0) := (others => '0');
    variable r2781 : std_logic_vector(0 to 0) := (others => '0');
    variable r2780 : std_logic_vector(0 to 0) := (others => '0');
    variable r2779 : std_logic_vector(0 to 0) := (others => '0');
    variable r2778 : std_logic_vector(0 to 0) := (others => '0');
    variable r2777 : std_logic_vector(0 to 0) := (others => '0');
    variable r2776 : std_logic_vector(0 to 0) := (others => '0');
    variable r2775 : std_logic_vector(0 to 0) := (others => '0');
    variable r2774 : std_logic_vector(0 to 0) := (others => '0');
    variable r2773 : std_logic_vector(0 to 0) := (others => '0');
    variable r2772 : std_logic_vector(0 to 0) := (others => '0');
    variable r2771 : std_logic_vector(0 to 0) := (others => '0');
    variable r2770 : std_logic_vector(0 to 0) := (others => '0');
    variable r2769 : std_logic_vector(0 to 0) := (others => '0');
    variable b2768 : boolean := false;
    variable r2767 : std_logic_vector(0 to 15) := (others => '0');
    variable r2766 : std_logic_vector(0 to 15) := (others => '0');
    variable b2765 : boolean := false;
    variable r2764 : std_logic_vector(0 to 31) := (others => '0');
    variable r2763 : std_logic_vector(0 to 31) := (others => '0');
  begin
    b2765 := true;
    r2766 := r2763(0 to 15);
    r2767 := r2763(16 to 31);
    b2768 := true;
    r2769 := r2766(0 to 0);
    r2770 := r2766(1 to 1);
    r2771 := r2766(2 to 2);
    r2772 := r2766(3 to 3);
    r2773 := r2766(4 to 4);
    r2774 := r2766(5 to 5);
    r2775 := r2766(6 to 6);
    r2776 := r2766(7 to 7);
    r2777 := r2766(8 to 8);
    r2778 := r2766(9 to 9);
    r2779 := r2766(10 to 10);
    r2780 := r2766(11 to 11);
    r2781 := r2766(12 to 12);
    r2782 := r2766(13 to 13);
    r2783 := r2766(14 to 14);
    r2784 := r2766(15 to 15);
    b2785 := true;
    b2786 := true;
    b2787 := true;
    b2788 := true;
    b2789 := true;
    b2790 := true;
    b2791 := true;
    b2792 := true;
    b2793 := true;
    b2794 := true;
    b2795 := true;
    b2796 := true;
    b2797 := true;
    b2798 := true;
    b2799 := true;
    b2800 := true;
    b2801 := (b2785 AND (b2786 AND (b2787 AND (b2788 AND (b2789 AND (b2790 AND (b2791 AND (b2792 AND (b2793 AND (b2794 AND (b2795 AND (b2796 AND (b2797 AND (b2798 AND (b2799 AND b2800)))))))))))))));
    b2802 := true;
    r2803 := r2767(0 to 0);
    r2804 := r2767(1 to 1);
    r2805 := r2767(2 to 2);
    r2806 := r2767(3 to 3);
    r2807 := r2767(4 to 4);
    r2808 := r2767(5 to 5);
    r2809 := r2767(6 to 6);
    r2810 := r2767(7 to 7);
    r2811 := r2767(8 to 8);
    r2812 := r2767(9 to 9);
    r2813 := r2767(10 to 10);
    r2814 := r2767(11 to 11);
    r2815 := r2767(12 to 12);
    r2816 := r2767(13 to 13);
    r2817 := r2767(14 to 14);
    r2818 := r2767(15 to 15);
    b2819 := true;
    b2820 := true;
    b2821 := true;
    b2822 := true;
    b2823 := true;
    b2824 := true;
    b2825 := true;
    b2826 := true;
    b2827 := true;
    b2828 := true;
    b2829 := true;
    b2830 := true;
    b2831 := true;
    b2832 := true;
    b2833 := true;
    b2834 := true;
    b2835 := (b2819 AND (b2820 AND (b2821 AND (b2822 AND (b2823 AND (b2824 AND (b2825 AND (b2826 AND (b2827 AND (b2828 AND (b2829 AND (b2830 AND (b2831 AND (b2832 AND (b2833 AND b2834)))))))))))))));
    b2836 := (b2801 AND b2835);
    if b2836 then
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      r2838 := (r2769 & r2770 & r2771 & r2772 & r2773 & r2774 & r2775 & r2776 & r2777 & r2778 & r2779 & r2780 & r2781 & r2782 & r2783 & r2784 & r2803 & r2804 & r2805 & r2806 & r2807 & r2808 & r2809 & r2810 & r2811 & r2812 & r2813 & r2814 & r2815 & r2816 & r2817 & r2818);
      r2764 := r2838;
    end if;
    return r2764;
  end rewire_w16tow32le_2758;
  function rewire_salsaHashp_1986(r1987 : std_logic_vector) return std_logic_vector
  is
    variable r2609 : std_logic_vector(0 to 511) := (others => '0');
    variable r2608 : std_logic_vector(0 to 31) := (others => '0');
    variable r2607 : std_logic_vector(0 to 31) := (others => '0');
    variable r2606 : std_logic_vector(0 to 31) := (others => '0');
    variable r2605 : std_logic_vector(0 to 31) := (others => '0');
    variable r2604 : std_logic_vector(0 to 31) := (others => '0');
    variable r2603 : std_logic_vector(0 to 31) := (others => '0');
    variable r2602 : std_logic_vector(0 to 31) := (others => '0');
    variable r2601 : std_logic_vector(0 to 31) := (others => '0');
    variable r2600 : std_logic_vector(0 to 31) := (others => '0');
    variable r2599 : std_logic_vector(0 to 31) := (others => '0');
    variable r2598 : std_logic_vector(0 to 31) := (others => '0');
    variable r2597 : std_logic_vector(0 to 31) := (others => '0');
    variable r2596 : std_logic_vector(0 to 31) := (others => '0');
    variable r2595 : std_logic_vector(0 to 31) := (others => '0');
    variable r2594 : std_logic_vector(0 to 31) := (others => '0');
    variable r2593 : std_logic_vector(0 to 31) := (others => '0');
    variable b2591 : boolean := false;
    variable b2590 : boolean := false;
    variable b2589 : boolean := false;
    variable b2588 : boolean := false;
    variable b2587 : boolean := false;
    variable b2586 : boolean := false;
    variable b2585 : boolean := false;
    variable b2584 : boolean := false;
    variable b2583 : boolean := false;
    variable b2582 : boolean := false;
    variable b2581 : boolean := false;
    variable b2580 : boolean := false;
    variable b2579 : boolean := false;
    variable b2578 : boolean := false;
    variable b2577 : boolean := false;
    variable b2576 : boolean := false;
    variable b2575 : boolean := false;
    variable r2574 : std_logic_vector(0 to 31) := (others => '0');
    variable r2573 : std_logic_vector(0 to 31) := (others => '0');
    variable r2572 : std_logic_vector(0 to 31) := (others => '0');
    variable r2571 : std_logic_vector(0 to 31) := (others => '0');
    variable r2570 : std_logic_vector(0 to 31) := (others => '0');
    variable r2569 : std_logic_vector(0 to 31) := (others => '0');
    variable r2568 : std_logic_vector(0 to 31) := (others => '0');
    variable r2567 : std_logic_vector(0 to 31) := (others => '0');
    variable r2566 : std_logic_vector(0 to 31) := (others => '0');
    variable r2565 : std_logic_vector(0 to 31) := (others => '0');
    variable r2564 : std_logic_vector(0 to 31) := (others => '0');
    variable r2563 : std_logic_vector(0 to 31) := (others => '0');
    variable r2562 : std_logic_vector(0 to 31) := (others => '0');
    variable r2561 : std_logic_vector(0 to 31) := (others => '0');
    variable r2560 : std_logic_vector(0 to 31) := (others => '0');
    variable r2559 : std_logic_vector(0 to 31) := (others => '0');
    variable b2558 : boolean := false;
    variable r2557 : std_logic_vector(0 to 511) := (others => '0');
    variable r2556 : std_logic_vector(0 to 511) := (others => '0');
    variable r2555 : std_logic_vector(0 to 511) := (others => '0');
    variable r2554 : std_logic_vector(0 to 511) := (others => '0');
    variable r2553 : std_logic_vector(0 to 511) := (others => '0');
    variable r2552 : std_logic_vector(0 to 511) := (others => '0');
    variable r2551 : std_logic_vector(0 to 511) := (others => '0');
    variable r2550 : std_logic_vector(0 to 511) := (others => '0');
    variable r2549 : std_logic_vector(0 to 511) := (others => '0');
    variable r2548 : std_logic_vector(0 to 511) := (others => '0');
    variable r2547 : std_logic_vector(0 to 511) := (others => '0');
    variable r2026 : std_logic_vector(0 to 511) := (others => '0');
    variable r2025 : std_logic_vector(0 to 511) := (others => '0');
    variable b2023 : boolean := false;
    variable b2022 : boolean := false;
    variable b2021 : boolean := false;
    variable b2020 : boolean := false;
    variable b2019 : boolean := false;
    variable b2018 : boolean := false;
    variable b2017 : boolean := false;
    variable b2016 : boolean := false;
    variable b2015 : boolean := false;
    variable b2014 : boolean := false;
    variable b2013 : boolean := false;
    variable b2012 : boolean := false;
    variable b2011 : boolean := false;
    variable b2010 : boolean := false;
    variable b2009 : boolean := false;
    variable b2008 : boolean := false;
    variable b2007 : boolean := false;
    variable r2006 : std_logic_vector(0 to 31) := (others => '0');
    variable r2005 : std_logic_vector(0 to 31) := (others => '0');
    variable r2004 : std_logic_vector(0 to 31) := (others => '0');
    variable r2003 : std_logic_vector(0 to 31) := (others => '0');
    variable r2002 : std_logic_vector(0 to 31) := (others => '0');
    variable r2001 : std_logic_vector(0 to 31) := (others => '0');
    variable r2000 : std_logic_vector(0 to 31) := (others => '0');
    variable r1999 : std_logic_vector(0 to 31) := (others => '0');
    variable r1998 : std_logic_vector(0 to 31) := (others => '0');
    variable r1997 : std_logic_vector(0 to 31) := (others => '0');
    variable r1996 : std_logic_vector(0 to 31) := (others => '0');
    variable r1995 : std_logic_vector(0 to 31) := (others => '0');
    variable r1994 : std_logic_vector(0 to 31) := (others => '0');
    variable r1993 : std_logic_vector(0 to 31) := (others => '0');
    variable r1992 : std_logic_vector(0 to 31) := (others => '0');
    variable r1991 : std_logic_vector(0 to 31) := (others => '0');
    variable b1990 : boolean := false;
    variable r1989 : std_logic_vector(0 to 511) := (others => '0');
  begin
    b1990 := true;
    r1991 := r1987(0 to 31);
    r1992 := r1987(32 to 63);
    r1993 := r1987(64 to 95);
    r1994 := r1987(96 to 127);
    r1995 := r1987(128 to 159);
    r1996 := r1987(160 to 191);
    r1997 := r1987(192 to 223);
    r1998 := r1987(224 to 255);
    r1999 := r1987(256 to 287);
    r2000 := r1987(288 to 319);
    r2001 := r1987(320 to 351);
    r2002 := r1987(352 to 383);
    r2003 := r1987(384 to 415);
    r2004 := r1987(416 to 447);
    r2005 := r1987(448 to 479);
    r2006 := r1987(480 to 511);
    b2007 := true;
    b2008 := true;
    b2009 := true;
    b2010 := true;
    b2011 := true;
    b2012 := true;
    b2013 := true;
    b2014 := true;
    b2015 := true;
    b2016 := true;
    b2017 := true;
    b2018 := true;
    b2019 := true;
    b2020 := true;
    b2021 := true;
    b2022 := true;
    b2023 := (b2007 AND (b2008 AND (b2009 AND (b2010 AND (b2011 AND (b2012 AND (b2013 AND (b2014 AND (b2015 AND (b2016 AND (b2017 AND (b2018 AND (b2019 AND (b2020 AND (b2021 AND b2022)))))))))))))));
    if b2023 then
      b2558 := true;
      r2559 := r2556(0 to 31);
      r2560 := r2556(32 to 63);
      r2561 := r2556(64 to 95);
      r2562 := r2556(96 to 127);
      r2563 := r2556(128 to 159);
      r2564 := r2556(160 to 191);
      r2565 := r2556(192 to 223);
      r2566 := r2556(224 to 255);
      r2567 := r2556(256 to 287);
      r2568 := r2556(288 to 319);
      r2569 := r2556(320 to 351);
      r2570 := r2556(352 to 383);
      r2571 := r2556(384 to 415);
      r2572 := r2556(416 to 447);
      r2573 := r2556(448 to 479);
      r2574 := r2556(480 to 511);
      b2575 := true;
      b2576 := true;
      b2577 := true;
      b2578 := true;
      b2579 := true;
      b2580 := true;
      b2581 := true;
      b2582 := true;
      b2583 := true;
      b2584 := true;
      b2585 := true;
      b2586 := true;
      b2587 := true;
      b2588 := true;
      b2589 := true;
      b2590 := true;
      b2591 := (b2575 AND (b2576 AND (b2577 AND (b2578 AND (b2579 AND (b2580 AND (b2581 AND (b2582 AND (b2583 AND (b2584 AND (b2585 AND (b2586 AND (b2587 AND (b2588 AND (b2589 AND b2590)))))))))))))));
      if b2591 then
        null;
        null;
        r2593 := add32(r2559,r1991);
        null;
        null;
        r2594 := add32(r2560,r1992);
        null;
        null;
        r2595 := add32(r2561,r1993);
        null;
        null;
        r2596 := add32(r2562,r1994);
        null;
        null;
        r2597 := add32(r2563,r1995);
        null;
        null;
        r2598 := add32(r2564,r1996);
        null;
        null;
        r2599 := add32(r2565,r1997);
        null;
        null;
        r2600 := add32(r2566,r1998);
        null;
        null;
        r2601 := add32(r2567,r1999);
        null;
        null;
        r2602 := add32(r2568,r2000);
        null;
        null;
        r2603 := add32(r2569,r2001);
        null;
        null;
        r2604 := add32(r2570,r2002);
        null;
        null;
        r2605 := add32(r2571,r2003);
        null;
        null;
        r2606 := add32(r2572,r2004);
        null;
        null;
        r2607 := add32(r2573,r2005);
        null;
        null;
        r2608 := add32(r2574,r2006);
        r2609 := (r2593 & r2594 & r2595 & r2596 & r2597 & r2598 & r2599 & r2600 & r2601 & r2602 & r2603 & r2604 & r2605 & r2606 & r2607 & r2608);
        r2557 := r2609;
      end if;
      r1989 := r2557;
    end if;
    return r1989;
  end rewire_salsaHashp_1986;
  function rewire_doubleRound_2024(r2025 : std_logic_vector) return std_logic_vector
  is
    variable r2546 : std_logic_vector(0 to 511) := (others => '0');
    variable r2545 : std_logic_vector(0 to 511) := (others => '0');
    variable r2446 : std_logic_vector(0 to 511) := (others => '0');
    variable r2445 : std_logic_vector(0 to 511) := (others => '0');
    variable r2029 : std_logic_vector(0 to 511) := (others => '0');
    variable r2028 : std_logic_vector(0 to 511) := (others => '0');
  begin
    null;
    r2545 := rewire_columnRound_2444(r2025);
    r2546 := rewire_rowRound_2027(r2545);
    return r2546;
  end rewire_doubleRound_2024;
  function rewire_columnRound_2444(r2445 : std_logic_vector) return std_logic_vector
  is
    variable r2544 : std_logic_vector(0 to 511) := (others => '0');
    variable b2542 : boolean := false;
    variable b2541 : boolean := false;
    variable b2540 : boolean := false;
    variable b2539 : boolean := false;
    variable b2538 : boolean := false;
    variable b2537 : boolean := false;
    variable r2536 : std_logic_vector(0 to 31) := (others => '0');
    variable r2535 : std_logic_vector(0 to 31) := (others => '0');
    variable r2534 : std_logic_vector(0 to 31) := (others => '0');
    variable r2533 : std_logic_vector(0 to 31) := (others => '0');
    variable b2532 : boolean := false;
    variable b2531 : boolean := false;
    variable b2530 : boolean := false;
    variable b2529 : boolean := false;
    variable b2528 : boolean := false;
    variable b2527 : boolean := false;
    variable r2526 : std_logic_vector(0 to 31) := (others => '0');
    variable r2525 : std_logic_vector(0 to 31) := (others => '0');
    variable r2524 : std_logic_vector(0 to 31) := (others => '0');
    variable r2523 : std_logic_vector(0 to 31) := (others => '0');
    variable b2522 : boolean := false;
    variable b2521 : boolean := false;
    variable b2520 : boolean := false;
    variable b2519 : boolean := false;
    variable b2518 : boolean := false;
    variable b2517 : boolean := false;
    variable r2516 : std_logic_vector(0 to 31) := (others => '0');
    variable r2515 : std_logic_vector(0 to 31) := (others => '0');
    variable r2514 : std_logic_vector(0 to 31) := (others => '0');
    variable r2513 : std_logic_vector(0 to 31) := (others => '0');
    variable b2512 : boolean := false;
    variable b2511 : boolean := false;
    variable b2510 : boolean := false;
    variable b2509 : boolean := false;
    variable b2508 : boolean := false;
    variable b2507 : boolean := false;
    variable r2506 : std_logic_vector(0 to 31) := (others => '0');
    variable r2505 : std_logic_vector(0 to 31) := (others => '0');
    variable r2504 : std_logic_vector(0 to 31) := (others => '0');
    variable r2503 : std_logic_vector(0 to 31) := (others => '0');
    variable b2502 : boolean := false;
    variable r2501 : std_logic_vector(0 to 127) := (others => '0');
    variable r2500 : std_logic_vector(0 to 127) := (others => '0');
    variable r2499 : std_logic_vector(0 to 127) := (others => '0');
    variable r2498 : std_logic_vector(0 to 127) := (others => '0');
    variable b2497 : boolean := false;
    variable r2496 : std_logic_vector(0 to 511) := (others => '0');
    variable r2495 : std_logic_vector(0 to 511) := (others => '0');
    variable r2493 : std_logic_vector(0 to 127) := (others => '0');
    variable r2492 : std_logic_vector(0 to 127) := (others => '0');
    variable r2490 : std_logic_vector(0 to 127) := (others => '0');
    variable r2489 : std_logic_vector(0 to 127) := (others => '0');
    variable r2487 : std_logic_vector(0 to 127) := (others => '0');
    variable r2486 : std_logic_vector(0 to 127) := (others => '0');
    variable r2484 : std_logic_vector(0 to 127) := (others => '0');
    variable r2483 : std_logic_vector(0 to 127) := (others => '0');
    variable b2481 : boolean := false;
    variable b2480 : boolean := false;
    variable b2479 : boolean := false;
    variable b2478 : boolean := false;
    variable b2477 : boolean := false;
    variable b2476 : boolean := false;
    variable b2475 : boolean := false;
    variable b2474 : boolean := false;
    variable b2473 : boolean := false;
    variable b2472 : boolean := false;
    variable b2471 : boolean := false;
    variable b2470 : boolean := false;
    variable b2469 : boolean := false;
    variable b2468 : boolean := false;
    variable b2467 : boolean := false;
    variable b2466 : boolean := false;
    variable b2465 : boolean := false;
    variable r2464 : std_logic_vector(0 to 31) := (others => '0');
    variable r2463 : std_logic_vector(0 to 31) := (others => '0');
    variable r2462 : std_logic_vector(0 to 31) := (others => '0');
    variable r2461 : std_logic_vector(0 to 31) := (others => '0');
    variable r2460 : std_logic_vector(0 to 31) := (others => '0');
    variable r2459 : std_logic_vector(0 to 31) := (others => '0');
    variable r2458 : std_logic_vector(0 to 31) := (others => '0');
    variable r2457 : std_logic_vector(0 to 31) := (others => '0');
    variable r2456 : std_logic_vector(0 to 31) := (others => '0');
    variable r2455 : std_logic_vector(0 to 31) := (others => '0');
    variable r2454 : std_logic_vector(0 to 31) := (others => '0');
    variable r2453 : std_logic_vector(0 to 31) := (others => '0');
    variable r2452 : std_logic_vector(0 to 31) := (others => '0');
    variable r2451 : std_logic_vector(0 to 31) := (others => '0');
    variable r2450 : std_logic_vector(0 to 31) := (others => '0');
    variable r2449 : std_logic_vector(0 to 31) := (others => '0');
    variable b2448 : boolean := false;
    variable r2447 : std_logic_vector(0 to 511) := (others => '0');
  begin
    b2448 := true;
    r2449 := r2445(0 to 31);
    r2450 := r2445(32 to 63);
    r2451 := r2445(64 to 95);
    r2452 := r2445(96 to 127);
    r2453 := r2445(128 to 159);
    r2454 := r2445(160 to 191);
    r2455 := r2445(192 to 223);
    r2456 := r2445(224 to 255);
    r2457 := r2445(256 to 287);
    r2458 := r2445(288 to 319);
    r2459 := r2445(320 to 351);
    r2460 := r2445(352 to 383);
    r2461 := r2445(384 to 415);
    r2462 := r2445(416 to 447);
    r2463 := r2445(448 to 479);
    r2464 := r2445(480 to 511);
    b2465 := true;
    b2466 := true;
    b2467 := true;
    b2468 := true;
    b2469 := true;
    b2470 := true;
    b2471 := true;
    b2472 := true;
    b2473 := true;
    b2474 := true;
    b2475 := true;
    b2476 := true;
    b2477 := true;
    b2478 := true;
    b2479 := true;
    b2480 := true;
    b2481 := (b2465 AND (b2466 AND (b2467 AND (b2468 AND (b2469 AND (b2470 AND (b2471 AND (b2472 AND (b2473 AND (b2474 AND (b2475 AND (b2476 AND (b2477 AND (b2478 AND (b2479 AND b2480)))))))))))))));
    if b2481 then
      null;
      null;
      null;
      null;
      r2483 := (r2449 & r2453 & r2457 & r2461);
      r2484 := rewire_quarterRound_2065(r2483);
      null;
      null;
      null;
      null;
      r2486 := (r2454 & r2458 & r2462 & r2450);
      r2487 := rewire_quarterRound_2065(r2486);
      null;
      null;
      null;
      null;
      r2489 := (r2459 & r2463 & r2451 & r2455);
      r2490 := rewire_quarterRound_2065(r2489);
      null;
      null;
      null;
      null;
      r2492 := (r2464 & r2452 & r2456 & r2460);
      r2493 := rewire_quarterRound_2065(r2492);
      b2497 := true;
      r2498 := r2495(0 to 127);
      r2499 := r2495(128 to 255);
      r2500 := r2495(256 to 383);
      r2501 := r2495(384 to 511);
      b2502 := true;
      r2503 := r2498(0 to 31);
      r2504 := r2498(32 to 63);
      r2505 := r2498(64 to 95);
      r2506 := r2498(96 to 127);
      b2507 := true;
      b2508 := true;
      b2509 := true;
      b2510 := true;
      b2511 := (b2507 AND (b2508 AND (b2509 AND b2510)));
      b2512 := true;
      r2513 := r2499(0 to 31);
      r2514 := r2499(32 to 63);
      r2515 := r2499(64 to 95);
      r2516 := r2499(96 to 127);
      b2517 := true;
      b2518 := true;
      b2519 := true;
      b2520 := true;
      b2521 := (b2517 AND (b2518 AND (b2519 AND b2520)));
      b2522 := true;
      r2523 := r2500(0 to 31);
      r2524 := r2500(32 to 63);
      r2525 := r2500(64 to 95);
      r2526 := r2500(96 to 127);
      b2527 := true;
      b2528 := true;
      b2529 := true;
      b2530 := true;
      b2531 := (b2527 AND (b2528 AND (b2529 AND b2530)));
      b2532 := true;
      r2533 := r2501(0 to 31);
      r2534 := r2501(32 to 63);
      r2535 := r2501(64 to 95);
      r2536 := r2501(96 to 127);
      b2537 := true;
      b2538 := true;
      b2539 := true;
      b2540 := true;
      b2541 := (b2537 AND (b2538 AND (b2539 AND b2540)));
      b2542 := (b2511 AND (b2521 AND (b2531 AND b2541)));
      if b2542 then
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        r2544 := (r2503 & r2516 & r2525 & r2534 & r2504 & r2513 & r2526 & r2535 & r2505 & r2514 & r2523 & r2536 & r2506 & r2515 & r2524 & r2533);
        r2496 := r2544;
      end if;
      r2447 := r2496;
    end if;
    return r2447;
  end rewire_columnRound_2444;
  function rewire_rowRound_2027(r2028 : std_logic_vector) return std_logic_vector
  is
    variable r2443 : std_logic_vector(0 to 511) := (others => '0');
    variable b2441 : boolean := false;
    variable b2440 : boolean := false;
    variable b2439 : boolean := false;
    variable b2438 : boolean := false;
    variable b2437 : boolean := false;
    variable b2436 : boolean := false;
    variable r2435 : std_logic_vector(0 to 31) := (others => '0');
    variable r2434 : std_logic_vector(0 to 31) := (others => '0');
    variable r2433 : std_logic_vector(0 to 31) := (others => '0');
    variable r2432 : std_logic_vector(0 to 31) := (others => '0');
    variable b2431 : boolean := false;
    variable b2430 : boolean := false;
    variable b2429 : boolean := false;
    variable b2428 : boolean := false;
    variable b2427 : boolean := false;
    variable b2426 : boolean := false;
    variable r2425 : std_logic_vector(0 to 31) := (others => '0');
    variable r2424 : std_logic_vector(0 to 31) := (others => '0');
    variable r2423 : std_logic_vector(0 to 31) := (others => '0');
    variable r2422 : std_logic_vector(0 to 31) := (others => '0');
    variable b2421 : boolean := false;
    variable b2420 : boolean := false;
    variable b2419 : boolean := false;
    variable b2418 : boolean := false;
    variable b2417 : boolean := false;
    variable b2416 : boolean := false;
    variable r2415 : std_logic_vector(0 to 31) := (others => '0');
    variable r2414 : std_logic_vector(0 to 31) := (others => '0');
    variable r2413 : std_logic_vector(0 to 31) := (others => '0');
    variable r2412 : std_logic_vector(0 to 31) := (others => '0');
    variable b2411 : boolean := false;
    variable b2410 : boolean := false;
    variable b2409 : boolean := false;
    variable b2408 : boolean := false;
    variable b2407 : boolean := false;
    variable b2406 : boolean := false;
    variable r2405 : std_logic_vector(0 to 31) := (others => '0');
    variable r2404 : std_logic_vector(0 to 31) := (others => '0');
    variable r2403 : std_logic_vector(0 to 31) := (others => '0');
    variable r2402 : std_logic_vector(0 to 31) := (others => '0');
    variable b2401 : boolean := false;
    variable r2400 : std_logic_vector(0 to 127) := (others => '0');
    variable r2399 : std_logic_vector(0 to 127) := (others => '0');
    variable r2398 : std_logic_vector(0 to 127) := (others => '0');
    variable r2397 : std_logic_vector(0 to 127) := (others => '0');
    variable b2396 : boolean := false;
    variable r2395 : std_logic_vector(0 to 511) := (others => '0');
    variable r2394 : std_logic_vector(0 to 511) := (others => '0');
    variable r2392 : std_logic_vector(0 to 127) := (others => '0');
    variable r2391 : std_logic_vector(0 to 127) := (others => '0');
    variable r2389 : std_logic_vector(0 to 127) := (others => '0');
    variable r2388 : std_logic_vector(0 to 127) := (others => '0');
    variable r2386 : std_logic_vector(0 to 127) := (others => '0');
    variable r2385 : std_logic_vector(0 to 127) := (others => '0');
    variable r2383 : std_logic_vector(0 to 127) := (others => '0');
    variable r2382 : std_logic_vector(0 to 127) := (others => '0');
    variable r2067 : std_logic_vector(0 to 127) := (others => '0');
    variable r2066 : std_logic_vector(0 to 127) := (others => '0');
    variable b2064 : boolean := false;
    variable b2063 : boolean := false;
    variable b2062 : boolean := false;
    variable b2061 : boolean := false;
    variable b2060 : boolean := false;
    variable b2059 : boolean := false;
    variable b2058 : boolean := false;
    variable b2057 : boolean := false;
    variable b2056 : boolean := false;
    variable b2055 : boolean := false;
    variable b2054 : boolean := false;
    variable b2053 : boolean := false;
    variable b2052 : boolean := false;
    variable b2051 : boolean := false;
    variable b2050 : boolean := false;
    variable b2049 : boolean := false;
    variable b2048 : boolean := false;
    variable r2047 : std_logic_vector(0 to 31) := (others => '0');
    variable r2046 : std_logic_vector(0 to 31) := (others => '0');
    variable r2045 : std_logic_vector(0 to 31) := (others => '0');
    variable r2044 : std_logic_vector(0 to 31) := (others => '0');
    variable r2043 : std_logic_vector(0 to 31) := (others => '0');
    variable r2042 : std_logic_vector(0 to 31) := (others => '0');
    variable r2041 : std_logic_vector(0 to 31) := (others => '0');
    variable r2040 : std_logic_vector(0 to 31) := (others => '0');
    variable r2039 : std_logic_vector(0 to 31) := (others => '0');
    variable r2038 : std_logic_vector(0 to 31) := (others => '0');
    variable r2037 : std_logic_vector(0 to 31) := (others => '0');
    variable r2036 : std_logic_vector(0 to 31) := (others => '0');
    variable r2035 : std_logic_vector(0 to 31) := (others => '0');
    variable r2034 : std_logic_vector(0 to 31) := (others => '0');
    variable r2033 : std_logic_vector(0 to 31) := (others => '0');
    variable r2032 : std_logic_vector(0 to 31) := (others => '0');
    variable b2031 : boolean := false;
    variable r2030 : std_logic_vector(0 to 511) := (others => '0');
  begin
    b2031 := true;
    r2032 := r2028(0 to 31);
    r2033 := r2028(32 to 63);
    r2034 := r2028(64 to 95);
    r2035 := r2028(96 to 127);
    r2036 := r2028(128 to 159);
    r2037 := r2028(160 to 191);
    r2038 := r2028(192 to 223);
    r2039 := r2028(224 to 255);
    r2040 := r2028(256 to 287);
    r2041 := r2028(288 to 319);
    r2042 := r2028(320 to 351);
    r2043 := r2028(352 to 383);
    r2044 := r2028(384 to 415);
    r2045 := r2028(416 to 447);
    r2046 := r2028(448 to 479);
    r2047 := r2028(480 to 511);
    b2048 := true;
    b2049 := true;
    b2050 := true;
    b2051 := true;
    b2052 := true;
    b2053 := true;
    b2054 := true;
    b2055 := true;
    b2056 := true;
    b2057 := true;
    b2058 := true;
    b2059 := true;
    b2060 := true;
    b2061 := true;
    b2062 := true;
    b2063 := true;
    b2064 := (b2048 AND (b2049 AND (b2050 AND (b2051 AND (b2052 AND (b2053 AND (b2054 AND (b2055 AND (b2056 AND (b2057 AND (b2058 AND (b2059 AND (b2060 AND (b2061 AND (b2062 AND b2063)))))))))))))));
    if b2064 then
      null;
      null;
      null;
      null;
      r2382 := (r2032 & r2033 & r2034 & r2035);
      r2383 := rewire_quarterRound_2065(r2382);
      null;
      null;
      null;
      null;
      r2385 := (r2037 & r2038 & r2039 & r2036);
      r2386 := rewire_quarterRound_2065(r2385);
      null;
      null;
      null;
      null;
      r2388 := (r2042 & r2043 & r2040 & r2041);
      r2389 := rewire_quarterRound_2065(r2388);
      null;
      null;
      null;
      null;
      r2391 := (r2047 & r2044 & r2045 & r2046);
      r2392 := rewire_quarterRound_2065(r2391);
      b2396 := true;
      r2397 := r2394(0 to 127);
      r2398 := r2394(128 to 255);
      r2399 := r2394(256 to 383);
      r2400 := r2394(384 to 511);
      b2401 := true;
      r2402 := r2397(0 to 31);
      r2403 := r2397(32 to 63);
      r2404 := r2397(64 to 95);
      r2405 := r2397(96 to 127);
      b2406 := true;
      b2407 := true;
      b2408 := true;
      b2409 := true;
      b2410 := (b2406 AND (b2407 AND (b2408 AND b2409)));
      b2411 := true;
      r2412 := r2398(0 to 31);
      r2413 := r2398(32 to 63);
      r2414 := r2398(64 to 95);
      r2415 := r2398(96 to 127);
      b2416 := true;
      b2417 := true;
      b2418 := true;
      b2419 := true;
      b2420 := (b2416 AND (b2417 AND (b2418 AND b2419)));
      b2421 := true;
      r2422 := r2399(0 to 31);
      r2423 := r2399(32 to 63);
      r2424 := r2399(64 to 95);
      r2425 := r2399(96 to 127);
      b2426 := true;
      b2427 := true;
      b2428 := true;
      b2429 := true;
      b2430 := (b2426 AND (b2427 AND (b2428 AND b2429)));
      b2431 := true;
      r2432 := r2400(0 to 31);
      r2433 := r2400(32 to 63);
      r2434 := r2400(64 to 95);
      r2435 := r2400(96 to 127);
      b2436 := true;
      b2437 := true;
      b2438 := true;
      b2439 := true;
      b2440 := (b2436 AND (b2437 AND (b2438 AND b2439)));
      b2441 := (b2410 AND (b2420 AND (b2430 AND b2440)));
      if b2441 then
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        r2443 := (r2402 & r2403 & r2404 & r2405 & r2415 & r2412 & r2413 & r2414 & r2424 & r2425 & r2422 & r2423 & r2433 & r2434 & r2435 & r2432);
        r2395 := r2443;
      end if;
      r2030 := r2395;
    end if;
    return r2030;
  end rewire_rowRound_2027;
  function rewire_quarterRound_2065(r2066 : std_logic_vector) return std_logic_vector
  is
    variable r2380 : std_logic_vector(0 to 127) := (others => '0');
    variable r2378 : std_logic_vector(0 to 31) := (others => '0');
    variable r2377 : std_logic_vector(0 to 31) := (others => '0');
    variable r2376 : std_logic_vector(0 to 31) := (others => '0');
    variable r2306 : std_logic_vector(0 to 31) := (others => '0');
    variable r2305 : std_logic_vector(0 to 31) := (others => '0');
    variable r2303 : std_logic_vector(0 to 31) := (others => '0');
    variable r2302 : std_logic_vector(0 to 31) := (others => '0');
    variable r2301 : std_logic_vector(0 to 31) := (others => '0');
    variable r2231 : std_logic_vector(0 to 31) := (others => '0');
    variable r2230 : std_logic_vector(0 to 31) := (others => '0');
    variable r2228 : std_logic_vector(0 to 31) := (others => '0');
    variable r2227 : std_logic_vector(0 to 31) := (others => '0');
    variable r2226 : std_logic_vector(0 to 31) := (others => '0');
    variable r2156 : std_logic_vector(0 to 31) := (others => '0');
    variable r2155 : std_logic_vector(0 to 31) := (others => '0');
    variable r2153 : std_logic_vector(0 to 31) := (others => '0');
    variable r2152 : std_logic_vector(0 to 31) := (others => '0');
    variable r2151 : std_logic_vector(0 to 31) := (others => '0');
    variable r2081 : std_logic_vector(0 to 31) := (others => '0');
    variable r2080 : std_logic_vector(0 to 31) := (others => '0');
    variable b2078 : boolean := false;
    variable b2077 : boolean := false;
    variable b2076 : boolean := false;
    variable b2075 : boolean := false;
    variable b2074 : boolean := false;
    variable r2073 : std_logic_vector(0 to 31) := (others => '0');
    variable r2072 : std_logic_vector(0 to 31) := (others => '0');
    variable r2071 : std_logic_vector(0 to 31) := (others => '0');
    variable r2070 : std_logic_vector(0 to 31) := (others => '0');
    variable b2069 : boolean := false;
    variable r2068 : std_logic_vector(0 to 127) := (others => '0');
  begin
    b2069 := true;
    r2070 := r2066(0 to 31);
    r2071 := r2066(32 to 63);
    r2072 := r2066(64 to 95);
    r2073 := r2066(96 to 127);
    b2074 := true;
    b2075 := true;
    b2076 := true;
    b2077 := true;
    b2078 := (b2074 AND (b2075 AND (b2076 AND b2077)));
    if b2078 then
      null;
      null;
      null;
      r2151 := add32(r2070,r2073);
      r2152 := rewire_rot7_2079(r2151);
      r2153 := xor32(r2071,r2152);
      null;
      null;
      null;
      r2226 := add32(r2153,r2070);
      r2227 := rewire_rot9_2154(r2226);
      r2228 := xor32(r2072,r2227);
      null;
      null;
      null;
      r2301 := add32(r2228,r2153);
      r2302 := rewire_rot13_2229(r2301);
      r2303 := xor32(r2073,r2302);
      null;
      null;
      null;
      r2376 := add32(r2303,r2228);
      r2377 := rewire_rot18_2304(r2376);
      r2378 := xor32(r2070,r2377);
      null;
      null;
      null;
      null;
      r2380 := (r2378 & r2153 & r2228 & r2303);
      r2068 := r2380;
    end if;
    return r2068;
  end rewire_quarterRound_2065;
  function rewire_rot18_2304(r2305 : std_logic_vector) return std_logic_vector
  is
    variable r2375 : std_logic_vector(0 to 31) := (others => '0');
    variable b2373 : boolean := false;
    variable b2372 : boolean := false;
    variable b2371 : boolean := false;
    variable b2370 : boolean := false;
    variable b2369 : boolean := false;
    variable b2368 : boolean := false;
    variable b2367 : boolean := false;
    variable b2366 : boolean := false;
    variable b2365 : boolean := false;
    variable b2364 : boolean := false;
    variable b2363 : boolean := false;
    variable b2362 : boolean := false;
    variable b2361 : boolean := false;
    variable b2360 : boolean := false;
    variable b2359 : boolean := false;
    variable b2358 : boolean := false;
    variable b2357 : boolean := false;
    variable b2356 : boolean := false;
    variable b2355 : boolean := false;
    variable b2354 : boolean := false;
    variable b2353 : boolean := false;
    variable b2352 : boolean := false;
    variable b2351 : boolean := false;
    variable b2350 : boolean := false;
    variable b2349 : boolean := false;
    variable b2348 : boolean := false;
    variable b2347 : boolean := false;
    variable b2346 : boolean := false;
    variable b2345 : boolean := false;
    variable b2344 : boolean := false;
    variable b2343 : boolean := false;
    variable b2342 : boolean := false;
    variable b2341 : boolean := false;
    variable r2340 : std_logic_vector(0 to 0) := (others => '0');
    variable r2339 : std_logic_vector(0 to 0) := (others => '0');
    variable r2338 : std_logic_vector(0 to 0) := (others => '0');
    variable r2337 : std_logic_vector(0 to 0) := (others => '0');
    variable r2336 : std_logic_vector(0 to 0) := (others => '0');
    variable r2335 : std_logic_vector(0 to 0) := (others => '0');
    variable r2334 : std_logic_vector(0 to 0) := (others => '0');
    variable r2333 : std_logic_vector(0 to 0) := (others => '0');
    variable r2332 : std_logic_vector(0 to 0) := (others => '0');
    variable r2331 : std_logic_vector(0 to 0) := (others => '0');
    variable r2330 : std_logic_vector(0 to 0) := (others => '0');
    variable r2329 : std_logic_vector(0 to 0) := (others => '0');
    variable r2328 : std_logic_vector(0 to 0) := (others => '0');
    variable r2327 : std_logic_vector(0 to 0) := (others => '0');
    variable r2326 : std_logic_vector(0 to 0) := (others => '0');
    variable r2325 : std_logic_vector(0 to 0) := (others => '0');
    variable r2324 : std_logic_vector(0 to 0) := (others => '0');
    variable r2323 : std_logic_vector(0 to 0) := (others => '0');
    variable r2322 : std_logic_vector(0 to 0) := (others => '0');
    variable r2321 : std_logic_vector(0 to 0) := (others => '0');
    variable r2320 : std_logic_vector(0 to 0) := (others => '0');
    variable r2319 : std_logic_vector(0 to 0) := (others => '0');
    variable r2318 : std_logic_vector(0 to 0) := (others => '0');
    variable r2317 : std_logic_vector(0 to 0) := (others => '0');
    variable r2316 : std_logic_vector(0 to 0) := (others => '0');
    variable r2315 : std_logic_vector(0 to 0) := (others => '0');
    variable r2314 : std_logic_vector(0 to 0) := (others => '0');
    variable r2313 : std_logic_vector(0 to 0) := (others => '0');
    variable r2312 : std_logic_vector(0 to 0) := (others => '0');
    variable r2311 : std_logic_vector(0 to 0) := (others => '0');
    variable r2310 : std_logic_vector(0 to 0) := (others => '0');
    variable r2309 : std_logic_vector(0 to 0) := (others => '0');
    variable b2308 : boolean := false;
    variable r2307 : std_logic_vector(0 to 31) := (others => '0');
  begin
    b2308 := true;
    r2309 := r2305(0 to 0);
    r2310 := r2305(1 to 1);
    r2311 := r2305(2 to 2);
    r2312 := r2305(3 to 3);
    r2313 := r2305(4 to 4);
    r2314 := r2305(5 to 5);
    r2315 := r2305(6 to 6);
    r2316 := r2305(7 to 7);
    r2317 := r2305(8 to 8);
    r2318 := r2305(9 to 9);
    r2319 := r2305(10 to 10);
    r2320 := r2305(11 to 11);
    r2321 := r2305(12 to 12);
    r2322 := r2305(13 to 13);
    r2323 := r2305(14 to 14);
    r2324 := r2305(15 to 15);
    r2325 := r2305(16 to 16);
    r2326 := r2305(17 to 17);
    r2327 := r2305(18 to 18);
    r2328 := r2305(19 to 19);
    r2329 := r2305(20 to 20);
    r2330 := r2305(21 to 21);
    r2331 := r2305(22 to 22);
    r2332 := r2305(23 to 23);
    r2333 := r2305(24 to 24);
    r2334 := r2305(25 to 25);
    r2335 := r2305(26 to 26);
    r2336 := r2305(27 to 27);
    r2337 := r2305(28 to 28);
    r2338 := r2305(29 to 29);
    r2339 := r2305(30 to 30);
    r2340 := r2305(31 to 31);
    b2341 := true;
    b2342 := true;
    b2343 := true;
    b2344 := true;
    b2345 := true;
    b2346 := true;
    b2347 := true;
    b2348 := true;
    b2349 := true;
    b2350 := true;
    b2351 := true;
    b2352 := true;
    b2353 := true;
    b2354 := true;
    b2355 := true;
    b2356 := true;
    b2357 := true;
    b2358 := true;
    b2359 := true;
    b2360 := true;
    b2361 := true;
    b2362 := true;
    b2363 := true;
    b2364 := true;
    b2365 := true;
    b2366 := true;
    b2367 := true;
    b2368 := true;
    b2369 := true;
    b2370 := true;
    b2371 := true;
    b2372 := true;
    b2373 := (b2341 AND (b2342 AND (b2343 AND (b2344 AND (b2345 AND (b2346 AND (b2347 AND (b2348 AND (b2349 AND (b2350 AND (b2351 AND (b2352 AND (b2353 AND (b2354 AND (b2355 AND (b2356 AND (b2357 AND (b2358 AND (b2359 AND (b2360 AND (b2361 AND (b2362 AND (b2363 AND (b2364 AND (b2365 AND (b2366 AND (b2367 AND (b2368 AND (b2369 AND (b2370 AND (b2371 AND b2372)))))))))))))))))))))))))))))));
    if b2373 then
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      r2375 := (r2327 & r2328 & r2329 & r2330 & r2331 & r2332 & r2333 & r2334 & r2335 & r2336 & r2337 & r2338 & r2339 & r2340 & r2309 & r2310 & r2311 & r2312 & r2313 & r2314 & r2315 & r2316 & r2317 & r2318 & r2319 & r2320 & r2321 & r2322 & r2323 & r2324 & r2325 & r2326);
      r2307 := r2375;
    end if;
    return r2307;
  end rewire_rot18_2304;
  function rewire_rot13_2229(r2230 : std_logic_vector) return std_logic_vector
  is
    variable r2300 : std_logic_vector(0 to 31) := (others => '0');
    variable b2298 : boolean := false;
    variable b2297 : boolean := false;
    variable b2296 : boolean := false;
    variable b2295 : boolean := false;
    variable b2294 : boolean := false;
    variable b2293 : boolean := false;
    variable b2292 : boolean := false;
    variable b2291 : boolean := false;
    variable b2290 : boolean := false;
    variable b2289 : boolean := false;
    variable b2288 : boolean := false;
    variable b2287 : boolean := false;
    variable b2286 : boolean := false;
    variable b2285 : boolean := false;
    variable b2284 : boolean := false;
    variable b2283 : boolean := false;
    variable b2282 : boolean := false;
    variable b2281 : boolean := false;
    variable b2280 : boolean := false;
    variable b2279 : boolean := false;
    variable b2278 : boolean := false;
    variable b2277 : boolean := false;
    variable b2276 : boolean := false;
    variable b2275 : boolean := false;
    variable b2274 : boolean := false;
    variable b2273 : boolean := false;
    variable b2272 : boolean := false;
    variable b2271 : boolean := false;
    variable b2270 : boolean := false;
    variable b2269 : boolean := false;
    variable b2268 : boolean := false;
    variable b2267 : boolean := false;
    variable b2266 : boolean := false;
    variable r2265 : std_logic_vector(0 to 0) := (others => '0');
    variable r2264 : std_logic_vector(0 to 0) := (others => '0');
    variable r2263 : std_logic_vector(0 to 0) := (others => '0');
    variable r2262 : std_logic_vector(0 to 0) := (others => '0');
    variable r2261 : std_logic_vector(0 to 0) := (others => '0');
    variable r2260 : std_logic_vector(0 to 0) := (others => '0');
    variable r2259 : std_logic_vector(0 to 0) := (others => '0');
    variable r2258 : std_logic_vector(0 to 0) := (others => '0');
    variable r2257 : std_logic_vector(0 to 0) := (others => '0');
    variable r2256 : std_logic_vector(0 to 0) := (others => '0');
    variable r2255 : std_logic_vector(0 to 0) := (others => '0');
    variable r2254 : std_logic_vector(0 to 0) := (others => '0');
    variable r2253 : std_logic_vector(0 to 0) := (others => '0');
    variable r2252 : std_logic_vector(0 to 0) := (others => '0');
    variable r2251 : std_logic_vector(0 to 0) := (others => '0');
    variable r2250 : std_logic_vector(0 to 0) := (others => '0');
    variable r2249 : std_logic_vector(0 to 0) := (others => '0');
    variable r2248 : std_logic_vector(0 to 0) := (others => '0');
    variable r2247 : std_logic_vector(0 to 0) := (others => '0');
    variable r2246 : std_logic_vector(0 to 0) := (others => '0');
    variable r2245 : std_logic_vector(0 to 0) := (others => '0');
    variable r2244 : std_logic_vector(0 to 0) := (others => '0');
    variable r2243 : std_logic_vector(0 to 0) := (others => '0');
    variable r2242 : std_logic_vector(0 to 0) := (others => '0');
    variable r2241 : std_logic_vector(0 to 0) := (others => '0');
    variable r2240 : std_logic_vector(0 to 0) := (others => '0');
    variable r2239 : std_logic_vector(0 to 0) := (others => '0');
    variable r2238 : std_logic_vector(0 to 0) := (others => '0');
    variable r2237 : std_logic_vector(0 to 0) := (others => '0');
    variable r2236 : std_logic_vector(0 to 0) := (others => '0');
    variable r2235 : std_logic_vector(0 to 0) := (others => '0');
    variable r2234 : std_logic_vector(0 to 0) := (others => '0');
    variable b2233 : boolean := false;
    variable r2232 : std_logic_vector(0 to 31) := (others => '0');
  begin
    b2233 := true;
    r2234 := r2230(0 to 0);
    r2235 := r2230(1 to 1);
    r2236 := r2230(2 to 2);
    r2237 := r2230(3 to 3);
    r2238 := r2230(4 to 4);
    r2239 := r2230(5 to 5);
    r2240 := r2230(6 to 6);
    r2241 := r2230(7 to 7);
    r2242 := r2230(8 to 8);
    r2243 := r2230(9 to 9);
    r2244 := r2230(10 to 10);
    r2245 := r2230(11 to 11);
    r2246 := r2230(12 to 12);
    r2247 := r2230(13 to 13);
    r2248 := r2230(14 to 14);
    r2249 := r2230(15 to 15);
    r2250 := r2230(16 to 16);
    r2251 := r2230(17 to 17);
    r2252 := r2230(18 to 18);
    r2253 := r2230(19 to 19);
    r2254 := r2230(20 to 20);
    r2255 := r2230(21 to 21);
    r2256 := r2230(22 to 22);
    r2257 := r2230(23 to 23);
    r2258 := r2230(24 to 24);
    r2259 := r2230(25 to 25);
    r2260 := r2230(26 to 26);
    r2261 := r2230(27 to 27);
    r2262 := r2230(28 to 28);
    r2263 := r2230(29 to 29);
    r2264 := r2230(30 to 30);
    r2265 := r2230(31 to 31);
    b2266 := true;
    b2267 := true;
    b2268 := true;
    b2269 := true;
    b2270 := true;
    b2271 := true;
    b2272 := true;
    b2273 := true;
    b2274 := true;
    b2275 := true;
    b2276 := true;
    b2277 := true;
    b2278 := true;
    b2279 := true;
    b2280 := true;
    b2281 := true;
    b2282 := true;
    b2283 := true;
    b2284 := true;
    b2285 := true;
    b2286 := true;
    b2287 := true;
    b2288 := true;
    b2289 := true;
    b2290 := true;
    b2291 := true;
    b2292 := true;
    b2293 := true;
    b2294 := true;
    b2295 := true;
    b2296 := true;
    b2297 := true;
    b2298 := (b2266 AND (b2267 AND (b2268 AND (b2269 AND (b2270 AND (b2271 AND (b2272 AND (b2273 AND (b2274 AND (b2275 AND (b2276 AND (b2277 AND (b2278 AND (b2279 AND (b2280 AND (b2281 AND (b2282 AND (b2283 AND (b2284 AND (b2285 AND (b2286 AND (b2287 AND (b2288 AND (b2289 AND (b2290 AND (b2291 AND (b2292 AND (b2293 AND (b2294 AND (b2295 AND (b2296 AND b2297)))))))))))))))))))))))))))))));
    if b2298 then
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      r2300 := (r2247 & r2248 & r2249 & r2250 & r2251 & r2252 & r2253 & r2254 & r2255 & r2256 & r2257 & r2258 & r2259 & r2260 & r2261 & r2262 & r2263 & r2264 & r2265 & r2234 & r2235 & r2236 & r2237 & r2238 & r2239 & r2240 & r2241 & r2242 & r2243 & r2244 & r2245 & r2246);
      r2232 := r2300;
    end if;
    return r2232;
  end rewire_rot13_2229;
  function rewire_rot9_2154(r2155 : std_logic_vector) return std_logic_vector
  is
    variable r2225 : std_logic_vector(0 to 31) := (others => '0');
    variable b2223 : boolean := false;
    variable b2222 : boolean := false;
    variable b2221 : boolean := false;
    variable b2220 : boolean := false;
    variable b2219 : boolean := false;
    variable b2218 : boolean := false;
    variable b2217 : boolean := false;
    variable b2216 : boolean := false;
    variable b2215 : boolean := false;
    variable b2214 : boolean := false;
    variable b2213 : boolean := false;
    variable b2212 : boolean := false;
    variable b2211 : boolean := false;
    variable b2210 : boolean := false;
    variable b2209 : boolean := false;
    variable b2208 : boolean := false;
    variable b2207 : boolean := false;
    variable b2206 : boolean := false;
    variable b2205 : boolean := false;
    variable b2204 : boolean := false;
    variable b2203 : boolean := false;
    variable b2202 : boolean := false;
    variable b2201 : boolean := false;
    variable b2200 : boolean := false;
    variable b2199 : boolean := false;
    variable b2198 : boolean := false;
    variable b2197 : boolean := false;
    variable b2196 : boolean := false;
    variable b2195 : boolean := false;
    variable b2194 : boolean := false;
    variable b2193 : boolean := false;
    variable b2192 : boolean := false;
    variable b2191 : boolean := false;
    variable r2190 : std_logic_vector(0 to 0) := (others => '0');
    variable r2189 : std_logic_vector(0 to 0) := (others => '0');
    variable r2188 : std_logic_vector(0 to 0) := (others => '0');
    variable r2187 : std_logic_vector(0 to 0) := (others => '0');
    variable r2186 : std_logic_vector(0 to 0) := (others => '0');
    variable r2185 : std_logic_vector(0 to 0) := (others => '0');
    variable r2184 : std_logic_vector(0 to 0) := (others => '0');
    variable r2183 : std_logic_vector(0 to 0) := (others => '0');
    variable r2182 : std_logic_vector(0 to 0) := (others => '0');
    variable r2181 : std_logic_vector(0 to 0) := (others => '0');
    variable r2180 : std_logic_vector(0 to 0) := (others => '0');
    variable r2179 : std_logic_vector(0 to 0) := (others => '0');
    variable r2178 : std_logic_vector(0 to 0) := (others => '0');
    variable r2177 : std_logic_vector(0 to 0) := (others => '0');
    variable r2176 : std_logic_vector(0 to 0) := (others => '0');
    variable r2175 : std_logic_vector(0 to 0) := (others => '0');
    variable r2174 : std_logic_vector(0 to 0) := (others => '0');
    variable r2173 : std_logic_vector(0 to 0) := (others => '0');
    variable r2172 : std_logic_vector(0 to 0) := (others => '0');
    variable r2171 : std_logic_vector(0 to 0) := (others => '0');
    variable r2170 : std_logic_vector(0 to 0) := (others => '0');
    variable r2169 : std_logic_vector(0 to 0) := (others => '0');
    variable r2168 : std_logic_vector(0 to 0) := (others => '0');
    variable r2167 : std_logic_vector(0 to 0) := (others => '0');
    variable r2166 : std_logic_vector(0 to 0) := (others => '0');
    variable r2165 : std_logic_vector(0 to 0) := (others => '0');
    variable r2164 : std_logic_vector(0 to 0) := (others => '0');
    variable r2163 : std_logic_vector(0 to 0) := (others => '0');
    variable r2162 : std_logic_vector(0 to 0) := (others => '0');
    variable r2161 : std_logic_vector(0 to 0) := (others => '0');
    variable r2160 : std_logic_vector(0 to 0) := (others => '0');
    variable r2159 : std_logic_vector(0 to 0) := (others => '0');
    variable b2158 : boolean := false;
    variable r2157 : std_logic_vector(0 to 31) := (others => '0');
  begin
    b2158 := true;
    r2159 := r2155(0 to 0);
    r2160 := r2155(1 to 1);
    r2161 := r2155(2 to 2);
    r2162 := r2155(3 to 3);
    r2163 := r2155(4 to 4);
    r2164 := r2155(5 to 5);
    r2165 := r2155(6 to 6);
    r2166 := r2155(7 to 7);
    r2167 := r2155(8 to 8);
    r2168 := r2155(9 to 9);
    r2169 := r2155(10 to 10);
    r2170 := r2155(11 to 11);
    r2171 := r2155(12 to 12);
    r2172 := r2155(13 to 13);
    r2173 := r2155(14 to 14);
    r2174 := r2155(15 to 15);
    r2175 := r2155(16 to 16);
    r2176 := r2155(17 to 17);
    r2177 := r2155(18 to 18);
    r2178 := r2155(19 to 19);
    r2179 := r2155(20 to 20);
    r2180 := r2155(21 to 21);
    r2181 := r2155(22 to 22);
    r2182 := r2155(23 to 23);
    r2183 := r2155(24 to 24);
    r2184 := r2155(25 to 25);
    r2185 := r2155(26 to 26);
    r2186 := r2155(27 to 27);
    r2187 := r2155(28 to 28);
    r2188 := r2155(29 to 29);
    r2189 := r2155(30 to 30);
    r2190 := r2155(31 to 31);
    b2191 := true;
    b2192 := true;
    b2193 := true;
    b2194 := true;
    b2195 := true;
    b2196 := true;
    b2197 := true;
    b2198 := true;
    b2199 := true;
    b2200 := true;
    b2201 := true;
    b2202 := true;
    b2203 := true;
    b2204 := true;
    b2205 := true;
    b2206 := true;
    b2207 := true;
    b2208 := true;
    b2209 := true;
    b2210 := true;
    b2211 := true;
    b2212 := true;
    b2213 := true;
    b2214 := true;
    b2215 := true;
    b2216 := true;
    b2217 := true;
    b2218 := true;
    b2219 := true;
    b2220 := true;
    b2221 := true;
    b2222 := true;
    b2223 := (b2191 AND (b2192 AND (b2193 AND (b2194 AND (b2195 AND (b2196 AND (b2197 AND (b2198 AND (b2199 AND (b2200 AND (b2201 AND (b2202 AND (b2203 AND (b2204 AND (b2205 AND (b2206 AND (b2207 AND (b2208 AND (b2209 AND (b2210 AND (b2211 AND (b2212 AND (b2213 AND (b2214 AND (b2215 AND (b2216 AND (b2217 AND (b2218 AND (b2219 AND (b2220 AND (b2221 AND b2222)))))))))))))))))))))))))))))));
    if b2223 then
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      r2225 := (r2168 & r2169 & r2170 & r2171 & r2172 & r2173 & r2174 & r2175 & r2176 & r2177 & r2178 & r2179 & r2180 & r2181 & r2182 & r2183 & r2184 & r2185 & r2186 & r2187 & r2188 & r2189 & r2190 & r2159 & r2160 & r2161 & r2162 & r2163 & r2164 & r2165 & r2166 & r2167);
      r2157 := r2225;
    end if;
    return r2157;
  end rewire_rot9_2154;
  function rewire_rot7_2079(r2080 : std_logic_vector) return std_logic_vector
  is
    variable r2150 : std_logic_vector(0 to 31) := (others => '0');
    variable b2148 : boolean := false;
    variable b2147 : boolean := false;
    variable b2146 : boolean := false;
    variable b2145 : boolean := false;
    variable b2144 : boolean := false;
    variable b2143 : boolean := false;
    variable b2142 : boolean := false;
    variable b2141 : boolean := false;
    variable b2140 : boolean := false;
    variable b2139 : boolean := false;
    variable b2138 : boolean := false;
    variable b2137 : boolean := false;
    variable b2136 : boolean := false;
    variable b2135 : boolean := false;
    variable b2134 : boolean := false;
    variable b2133 : boolean := false;
    variable b2132 : boolean := false;
    variable b2131 : boolean := false;
    variable b2130 : boolean := false;
    variable b2129 : boolean := false;
    variable b2128 : boolean := false;
    variable b2127 : boolean := false;
    variable b2126 : boolean := false;
    variable b2125 : boolean := false;
    variable b2124 : boolean := false;
    variable b2123 : boolean := false;
    variable b2122 : boolean := false;
    variable b2121 : boolean := false;
    variable b2120 : boolean := false;
    variable b2119 : boolean := false;
    variable b2118 : boolean := false;
    variable b2117 : boolean := false;
    variable b2116 : boolean := false;
    variable r2115 : std_logic_vector(0 to 0) := (others => '0');
    variable r2114 : std_logic_vector(0 to 0) := (others => '0');
    variable r2113 : std_logic_vector(0 to 0) := (others => '0');
    variable r2112 : std_logic_vector(0 to 0) := (others => '0');
    variable r2111 : std_logic_vector(0 to 0) := (others => '0');
    variable r2110 : std_logic_vector(0 to 0) := (others => '0');
    variable r2109 : std_logic_vector(0 to 0) := (others => '0');
    variable r2108 : std_logic_vector(0 to 0) := (others => '0');
    variable r2107 : std_logic_vector(0 to 0) := (others => '0');
    variable r2106 : std_logic_vector(0 to 0) := (others => '0');
    variable r2105 : std_logic_vector(0 to 0) := (others => '0');
    variable r2104 : std_logic_vector(0 to 0) := (others => '0');
    variable r2103 : std_logic_vector(0 to 0) := (others => '0');
    variable r2102 : std_logic_vector(0 to 0) := (others => '0');
    variable r2101 : std_logic_vector(0 to 0) := (others => '0');
    variable r2100 : std_logic_vector(0 to 0) := (others => '0');
    variable r2099 : std_logic_vector(0 to 0) := (others => '0');
    variable r2098 : std_logic_vector(0 to 0) := (others => '0');
    variable r2097 : std_logic_vector(0 to 0) := (others => '0');
    variable r2096 : std_logic_vector(0 to 0) := (others => '0');
    variable r2095 : std_logic_vector(0 to 0) := (others => '0');
    variable r2094 : std_logic_vector(0 to 0) := (others => '0');
    variable r2093 : std_logic_vector(0 to 0) := (others => '0');
    variable r2092 : std_logic_vector(0 to 0) := (others => '0');
    variable r2091 : std_logic_vector(0 to 0) := (others => '0');
    variable r2090 : std_logic_vector(0 to 0) := (others => '0');
    variable r2089 : std_logic_vector(0 to 0) := (others => '0');
    variable r2088 : std_logic_vector(0 to 0) := (others => '0');
    variable r2087 : std_logic_vector(0 to 0) := (others => '0');
    variable r2086 : std_logic_vector(0 to 0) := (others => '0');
    variable r2085 : std_logic_vector(0 to 0) := (others => '0');
    variable r2084 : std_logic_vector(0 to 0) := (others => '0');
    variable b2083 : boolean := false;
    variable r2082 : std_logic_vector(0 to 31) := (others => '0');
  begin
    b2083 := true;
    r2084 := r2080(0 to 0);
    r2085 := r2080(1 to 1);
    r2086 := r2080(2 to 2);
    r2087 := r2080(3 to 3);
    r2088 := r2080(4 to 4);
    r2089 := r2080(5 to 5);
    r2090 := r2080(6 to 6);
    r2091 := r2080(7 to 7);
    r2092 := r2080(8 to 8);
    r2093 := r2080(9 to 9);
    r2094 := r2080(10 to 10);
    r2095 := r2080(11 to 11);
    r2096 := r2080(12 to 12);
    r2097 := r2080(13 to 13);
    r2098 := r2080(14 to 14);
    r2099 := r2080(15 to 15);
    r2100 := r2080(16 to 16);
    r2101 := r2080(17 to 17);
    r2102 := r2080(18 to 18);
    r2103 := r2080(19 to 19);
    r2104 := r2080(20 to 20);
    r2105 := r2080(21 to 21);
    r2106 := r2080(22 to 22);
    r2107 := r2080(23 to 23);
    r2108 := r2080(24 to 24);
    r2109 := r2080(25 to 25);
    r2110 := r2080(26 to 26);
    r2111 := r2080(27 to 27);
    r2112 := r2080(28 to 28);
    r2113 := r2080(29 to 29);
    r2114 := r2080(30 to 30);
    r2115 := r2080(31 to 31);
    b2116 := true;
    b2117 := true;
    b2118 := true;
    b2119 := true;
    b2120 := true;
    b2121 := true;
    b2122 := true;
    b2123 := true;
    b2124 := true;
    b2125 := true;
    b2126 := true;
    b2127 := true;
    b2128 := true;
    b2129 := true;
    b2130 := true;
    b2131 := true;
    b2132 := true;
    b2133 := true;
    b2134 := true;
    b2135 := true;
    b2136 := true;
    b2137 := true;
    b2138 := true;
    b2139 := true;
    b2140 := true;
    b2141 := true;
    b2142 := true;
    b2143 := true;
    b2144 := true;
    b2145 := true;
    b2146 := true;
    b2147 := true;
    b2148 := (b2116 AND (b2117 AND (b2118 AND (b2119 AND (b2120 AND (b2121 AND (b2122 AND (b2123 AND (b2124 AND (b2125 AND (b2126 AND (b2127 AND (b2128 AND (b2129 AND (b2130 AND (b2131 AND (b2132 AND (b2133 AND (b2134 AND (b2135 AND (b2136 AND (b2137 AND (b2138 AND (b2139 AND (b2140 AND (b2141 AND (b2142 AND (b2143 AND (b2144 AND (b2145 AND (b2146 AND b2147)))))))))))))))))))))))))))))));
    if b2148 then
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      r2150 := (r2091 & r2092 & r2093 & r2094 & r2095 & r2096 & r2097 & r2098 & r2099 & r2100 & r2101 & r2102 & r2103 & r2104 & r2105 & r2106 & r2107 & r2108 & r2109 & r2110 & r2111 & r2112 & r2113 & r2114 & r2115 & r2084 & r2085 & r2086 & r2087 & r2088 & r2089 & r2090);
      r2082 := r2150;
    end if;
    return r2082;
  end rewire_rot7_2079;
  function rewire_expwords_1669(r1670 : std_logic_vector) return std_logic_vector
  is
    variable r1985 : std_logic_vector(0 to 511) := (others => '0');
    variable b1983 : boolean := false;
    variable b1982 : boolean := false;
    variable b1981 : boolean := false;
    variable b1980 : boolean := false;
    variable b1979 : boolean := false;
    variable b1978 : boolean := false;
    variable r1977 : std_logic_vector(0 to 7) := (others => '0');
    variable r1976 : std_logic_vector(0 to 7) := (others => '0');
    variable r1975 : std_logic_vector(0 to 7) := (others => '0');
    variable r1974 : std_logic_vector(0 to 7) := (others => '0');
    variable b1973 : boolean := false;
    variable b1972 : boolean := false;
    variable b1971 : boolean := false;
    variable b1970 : boolean := false;
    variable b1969 : boolean := false;
    variable b1968 : boolean := false;
    variable r1967 : std_logic_vector(0 to 7) := (others => '0');
    variable r1966 : std_logic_vector(0 to 7) := (others => '0');
    variable r1965 : std_logic_vector(0 to 7) := (others => '0');
    variable r1964 : std_logic_vector(0 to 7) := (others => '0');
    variable b1963 : boolean := false;
    variable b1962 : boolean := false;
    variable b1961 : boolean := false;
    variable b1960 : boolean := false;
    variable b1959 : boolean := false;
    variable b1958 : boolean := false;
    variable r1957 : std_logic_vector(0 to 7) := (others => '0');
    variable r1956 : std_logic_vector(0 to 7) := (others => '0');
    variable r1955 : std_logic_vector(0 to 7) := (others => '0');
    variable r1954 : std_logic_vector(0 to 7) := (others => '0');
    variable b1953 : boolean := false;
    variable b1952 : boolean := false;
    variable b1951 : boolean := false;
    variable b1950 : boolean := false;
    variable b1949 : boolean := false;
    variable b1948 : boolean := false;
    variable r1947 : std_logic_vector(0 to 7) := (others => '0');
    variable r1946 : std_logic_vector(0 to 7) := (others => '0');
    variable r1945 : std_logic_vector(0 to 7) := (others => '0');
    variable r1944 : std_logic_vector(0 to 7) := (others => '0');
    variable b1943 : boolean := false;
    variable b1942 : boolean := false;
    variable b1941 : boolean := false;
    variable b1940 : boolean := false;
    variable b1939 : boolean := false;
    variable b1938 : boolean := false;
    variable r1937 : std_logic_vector(0 to 7) := (others => '0');
    variable r1936 : std_logic_vector(0 to 7) := (others => '0');
    variable r1935 : std_logic_vector(0 to 7) := (others => '0');
    variable r1934 : std_logic_vector(0 to 7) := (others => '0');
    variable b1933 : boolean := false;
    variable b1932 : boolean := false;
    variable b1931 : boolean := false;
    variable b1930 : boolean := false;
    variable b1929 : boolean := false;
    variable b1928 : boolean := false;
    variable r1927 : std_logic_vector(0 to 7) := (others => '0');
    variable r1926 : std_logic_vector(0 to 7) := (others => '0');
    variable r1925 : std_logic_vector(0 to 7) := (others => '0');
    variable r1924 : std_logic_vector(0 to 7) := (others => '0');
    variable b1923 : boolean := false;
    variable b1922 : boolean := false;
    variable b1921 : boolean := false;
    variable b1920 : boolean := false;
    variable b1919 : boolean := false;
    variable b1918 : boolean := false;
    variable r1917 : std_logic_vector(0 to 7) := (others => '0');
    variable r1916 : std_logic_vector(0 to 7) := (others => '0');
    variable r1915 : std_logic_vector(0 to 7) := (others => '0');
    variable r1914 : std_logic_vector(0 to 7) := (others => '0');
    variable b1913 : boolean := false;
    variable b1912 : boolean := false;
    variable b1911 : boolean := false;
    variable b1910 : boolean := false;
    variable b1909 : boolean := false;
    variable b1908 : boolean := false;
    variable r1907 : std_logic_vector(0 to 7) := (others => '0');
    variable r1906 : std_logic_vector(0 to 7) := (others => '0');
    variable r1905 : std_logic_vector(0 to 7) := (others => '0');
    variable r1904 : std_logic_vector(0 to 7) := (others => '0');
    variable b1903 : boolean := false;
    variable b1902 : boolean := false;
    variable b1901 : boolean := false;
    variable b1900 : boolean := false;
    variable b1899 : boolean := false;
    variable b1898 : boolean := false;
    variable r1897 : std_logic_vector(0 to 7) := (others => '0');
    variable r1896 : std_logic_vector(0 to 7) := (others => '0');
    variable r1895 : std_logic_vector(0 to 7) := (others => '0');
    variable r1894 : std_logic_vector(0 to 7) := (others => '0');
    variable b1893 : boolean := false;
    variable b1892 : boolean := false;
    variable b1891 : boolean := false;
    variable b1890 : boolean := false;
    variable b1889 : boolean := false;
    variable b1888 : boolean := false;
    variable r1887 : std_logic_vector(0 to 7) := (others => '0');
    variable r1886 : std_logic_vector(0 to 7) := (others => '0');
    variable r1885 : std_logic_vector(0 to 7) := (others => '0');
    variable r1884 : std_logic_vector(0 to 7) := (others => '0');
    variable b1883 : boolean := false;
    variable b1882 : boolean := false;
    variable b1881 : boolean := false;
    variable b1880 : boolean := false;
    variable b1879 : boolean := false;
    variable b1878 : boolean := false;
    variable r1877 : std_logic_vector(0 to 7) := (others => '0');
    variable r1876 : std_logic_vector(0 to 7) := (others => '0');
    variable r1875 : std_logic_vector(0 to 7) := (others => '0');
    variable r1874 : std_logic_vector(0 to 7) := (others => '0');
    variable b1873 : boolean := false;
    variable b1872 : boolean := false;
    variable b1871 : boolean := false;
    variable b1870 : boolean := false;
    variable b1869 : boolean := false;
    variable b1868 : boolean := false;
    variable r1867 : std_logic_vector(0 to 7) := (others => '0');
    variable r1866 : std_logic_vector(0 to 7) := (others => '0');
    variable r1865 : std_logic_vector(0 to 7) := (others => '0');
    variable r1864 : std_logic_vector(0 to 7) := (others => '0');
    variable b1863 : boolean := false;
    variable b1862 : boolean := false;
    variable b1861 : boolean := false;
    variable b1860 : boolean := false;
    variable b1859 : boolean := false;
    variable b1858 : boolean := false;
    variable r1857 : std_logic_vector(0 to 7) := (others => '0');
    variable r1856 : std_logic_vector(0 to 7) := (others => '0');
    variable r1855 : std_logic_vector(0 to 7) := (others => '0');
    variable r1854 : std_logic_vector(0 to 7) := (others => '0');
    variable b1853 : boolean := false;
    variable b1852 : boolean := false;
    variable b1851 : boolean := false;
    variable b1850 : boolean := false;
    variable b1849 : boolean := false;
    variable b1848 : boolean := false;
    variable r1847 : std_logic_vector(0 to 7) := (others => '0');
    variable r1846 : std_logic_vector(0 to 7) := (others => '0');
    variable r1845 : std_logic_vector(0 to 7) := (others => '0');
    variable r1844 : std_logic_vector(0 to 7) := (others => '0');
    variable b1843 : boolean := false;
    variable b1842 : boolean := false;
    variable b1841 : boolean := false;
    variable b1840 : boolean := false;
    variable b1839 : boolean := false;
    variable b1838 : boolean := false;
    variable r1837 : std_logic_vector(0 to 7) := (others => '0');
    variable r1836 : std_logic_vector(0 to 7) := (others => '0');
    variable r1835 : std_logic_vector(0 to 7) := (others => '0');
    variable r1834 : std_logic_vector(0 to 7) := (others => '0');
    variable b1833 : boolean := false;
    variable b1832 : boolean := false;
    variable b1831 : boolean := false;
    variable b1830 : boolean := false;
    variable b1829 : boolean := false;
    variable b1828 : boolean := false;
    variable r1827 : std_logic_vector(0 to 7) := (others => '0');
    variable r1826 : std_logic_vector(0 to 7) := (others => '0');
    variable r1825 : std_logic_vector(0 to 7) := (others => '0');
    variable r1824 : std_logic_vector(0 to 7) := (others => '0');
    variable b1823 : boolean := false;
    variable r1822 : std_logic_vector(0 to 31) := (others => '0');
    variable r1821 : std_logic_vector(0 to 31) := (others => '0');
    variable r1820 : std_logic_vector(0 to 31) := (others => '0');
    variable r1819 : std_logic_vector(0 to 31) := (others => '0');
    variable r1818 : std_logic_vector(0 to 31) := (others => '0');
    variable r1817 : std_logic_vector(0 to 31) := (others => '0');
    variable r1816 : std_logic_vector(0 to 31) := (others => '0');
    variable r1815 : std_logic_vector(0 to 31) := (others => '0');
    variable r1814 : std_logic_vector(0 to 31) := (others => '0');
    variable r1813 : std_logic_vector(0 to 31) := (others => '0');
    variable r1812 : std_logic_vector(0 to 31) := (others => '0');
    variable r1811 : std_logic_vector(0 to 31) := (others => '0');
    variable r1810 : std_logic_vector(0 to 31) := (others => '0');
    variable r1809 : std_logic_vector(0 to 31) := (others => '0');
    variable r1808 : std_logic_vector(0 to 31) := (others => '0');
    variable r1807 : std_logic_vector(0 to 31) := (others => '0');
    variable b1806 : boolean := false;
    variable r1805 : std_logic_vector(0 to 511) := (others => '0');
    variable r1804 : std_logic_vector(0 to 511) := (others => '0');
    variable r1802 : std_logic_vector(0 to 31) := (others => '0');
    variable r1801 : std_logic_vector(0 to 31) := (others => '0');
    variable r1800 : std_logic_vector(0 to 31) := (others => '0');
    variable r1799 : std_logic_vector(0 to 31) := (others => '0');
    variable r1798 : std_logic_vector(0 to 31) := (others => '0');
    variable r1797 : std_logic_vector(0 to 31) := (others => '0');
    variable r1796 : std_logic_vector(0 to 31) := (others => '0');
    variable r1795 : std_logic_vector(0 to 31) := (others => '0');
    variable r1794 : std_logic_vector(0 to 31) := (others => '0');
    variable r1793 : std_logic_vector(0 to 31) := (others => '0');
    variable r1792 : std_logic_vector(0 to 31) := (others => '0');
    variable r1791 : std_logic_vector(0 to 31) := (others => '0');
    variable r1790 : std_logic_vector(0 to 31) := (others => '0');
    variable r1789 : std_logic_vector(0 to 31) := (others => '0');
    variable r1788 : std_logic_vector(0 to 31) := (others => '0');
    variable r1787 : std_logic_vector(0 to 31) := (others => '0');
    variable r1709 : std_logic_vector(0 to 31) := (others => '0');
    variable r1708 : std_logic_vector(0 to 31) := (others => '0');
    variable b1706 : boolean := false;
    variable b1705 : boolean := false;
    variable b1704 : boolean := false;
    variable b1703 : boolean := false;
    variable b1702 : boolean := false;
    variable b1701 : boolean := false;
    variable b1700 : boolean := false;
    variable b1699 : boolean := false;
    variable b1698 : boolean := false;
    variable b1697 : boolean := false;
    variable b1696 : boolean := false;
    variable b1695 : boolean := false;
    variable b1694 : boolean := false;
    variable b1693 : boolean := false;
    variable b1692 : boolean := false;
    variable b1691 : boolean := false;
    variable b1690 : boolean := false;
    variable r1689 : std_logic_vector(0 to 31) := (others => '0');
    variable r1688 : std_logic_vector(0 to 31) := (others => '0');
    variable r1687 : std_logic_vector(0 to 31) := (others => '0');
    variable r1686 : std_logic_vector(0 to 31) := (others => '0');
    variable r1685 : std_logic_vector(0 to 31) := (others => '0');
    variable r1684 : std_logic_vector(0 to 31) := (others => '0');
    variable r1683 : std_logic_vector(0 to 31) := (others => '0');
    variable r1682 : std_logic_vector(0 to 31) := (others => '0');
    variable r1681 : std_logic_vector(0 to 31) := (others => '0');
    variable r1680 : std_logic_vector(0 to 31) := (others => '0');
    variable r1679 : std_logic_vector(0 to 31) := (others => '0');
    variable r1678 : std_logic_vector(0 to 31) := (others => '0');
    variable r1677 : std_logic_vector(0 to 31) := (others => '0');
    variable r1676 : std_logic_vector(0 to 31) := (others => '0');
    variable r1675 : std_logic_vector(0 to 31) := (others => '0');
    variable r1674 : std_logic_vector(0 to 31) := (others => '0');
    variable b1673 : boolean := false;
    variable r1672 : std_logic_vector(0 to 511) := (others => '0');
  begin
    b1673 := true;
    r1674 := r1670(0 to 31);
    r1675 := r1670(32 to 63);
    r1676 := r1670(64 to 95);
    r1677 := r1670(96 to 127);
    r1678 := r1670(128 to 159);
    r1679 := r1670(160 to 191);
    r1680 := r1670(192 to 223);
    r1681 := r1670(224 to 255);
    r1682 := r1670(256 to 287);
    r1683 := r1670(288 to 319);
    r1684 := r1670(320 to 351);
    r1685 := r1670(352 to 383);
    r1686 := r1670(384 to 415);
    r1687 := r1670(416 to 447);
    r1688 := r1670(448 to 479);
    r1689 := r1670(480 to 511);
    b1690 := true;
    b1691 := true;
    b1692 := true;
    b1693 := true;
    b1694 := true;
    b1695 := true;
    b1696 := true;
    b1697 := true;
    b1698 := true;
    b1699 := true;
    b1700 := true;
    b1701 := true;
    b1702 := true;
    b1703 := true;
    b1704 := true;
    b1705 := true;
    b1706 := (b1690 AND (b1691 AND (b1692 AND (b1693 AND (b1694 AND (b1695 AND (b1696 AND (b1697 AND (b1698 AND (b1699 AND (b1700 AND (b1701 AND (b1702 AND (b1703 AND (b1704 AND b1705)))))))))))))));
    if b1706 then
      null;
      r1787 := rewire_littleendianp_1707(r1674);
      null;
      r1788 := rewire_littleendianp_1707(r1675);
      null;
      r1789 := rewire_littleendianp_1707(r1676);
      null;
      r1790 := rewire_littleendianp_1707(r1677);
      null;
      r1791 := rewire_littleendianp_1707(r1678);
      null;
      r1792 := rewire_littleendianp_1707(r1679);
      null;
      r1793 := rewire_littleendianp_1707(r1680);
      null;
      r1794 := rewire_littleendianp_1707(r1681);
      null;
      r1795 := rewire_littleendianp_1707(r1682);
      null;
      r1796 := rewire_littleendianp_1707(r1683);
      null;
      r1797 := rewire_littleendianp_1707(r1684);
      null;
      r1798 := rewire_littleendianp_1707(r1685);
      null;
      r1799 := rewire_littleendianp_1707(r1686);
      null;
      r1800 := rewire_littleendianp_1707(r1687);
      null;
      r1801 := rewire_littleendianp_1707(r1688);
      null;
      r1802 := rewire_littleendianp_1707(r1689);
      b1806 := true;
      r1807 := r1804(0 to 31);
      r1808 := r1804(32 to 63);
      r1809 := r1804(64 to 95);
      r1810 := r1804(96 to 127);
      r1811 := r1804(128 to 159);
      r1812 := r1804(160 to 191);
      r1813 := r1804(192 to 223);
      r1814 := r1804(224 to 255);
      r1815 := r1804(256 to 287);
      r1816 := r1804(288 to 319);
      r1817 := r1804(320 to 351);
      r1818 := r1804(352 to 383);
      r1819 := r1804(384 to 415);
      r1820 := r1804(416 to 447);
      r1821 := r1804(448 to 479);
      r1822 := r1804(480 to 511);
      b1823 := true;
      r1824 := r1807(0 to 7);
      r1825 := r1807(8 to 15);
      r1826 := r1807(16 to 23);
      r1827 := r1807(24 to 31);
      b1828 := true;
      b1829 := true;
      b1830 := true;
      b1831 := true;
      b1832 := (b1828 AND (b1829 AND (b1830 AND b1831)));
      b1833 := true;
      r1834 := r1808(0 to 7);
      r1835 := r1808(8 to 15);
      r1836 := r1808(16 to 23);
      r1837 := r1808(24 to 31);
      b1838 := true;
      b1839 := true;
      b1840 := true;
      b1841 := true;
      b1842 := (b1838 AND (b1839 AND (b1840 AND b1841)));
      b1843 := true;
      r1844 := r1809(0 to 7);
      r1845 := r1809(8 to 15);
      r1846 := r1809(16 to 23);
      r1847 := r1809(24 to 31);
      b1848 := true;
      b1849 := true;
      b1850 := true;
      b1851 := true;
      b1852 := (b1848 AND (b1849 AND (b1850 AND b1851)));
      b1853 := true;
      r1854 := r1810(0 to 7);
      r1855 := r1810(8 to 15);
      r1856 := r1810(16 to 23);
      r1857 := r1810(24 to 31);
      b1858 := true;
      b1859 := true;
      b1860 := true;
      b1861 := true;
      b1862 := (b1858 AND (b1859 AND (b1860 AND b1861)));
      b1863 := true;
      r1864 := r1811(0 to 7);
      r1865 := r1811(8 to 15);
      r1866 := r1811(16 to 23);
      r1867 := r1811(24 to 31);
      b1868 := true;
      b1869 := true;
      b1870 := true;
      b1871 := true;
      b1872 := (b1868 AND (b1869 AND (b1870 AND b1871)));
      b1873 := true;
      r1874 := r1812(0 to 7);
      r1875 := r1812(8 to 15);
      r1876 := r1812(16 to 23);
      r1877 := r1812(24 to 31);
      b1878 := true;
      b1879 := true;
      b1880 := true;
      b1881 := true;
      b1882 := (b1878 AND (b1879 AND (b1880 AND b1881)));
      b1883 := true;
      r1884 := r1813(0 to 7);
      r1885 := r1813(8 to 15);
      r1886 := r1813(16 to 23);
      r1887 := r1813(24 to 31);
      b1888 := true;
      b1889 := true;
      b1890 := true;
      b1891 := true;
      b1892 := (b1888 AND (b1889 AND (b1890 AND b1891)));
      b1893 := true;
      r1894 := r1814(0 to 7);
      r1895 := r1814(8 to 15);
      r1896 := r1814(16 to 23);
      r1897 := r1814(24 to 31);
      b1898 := true;
      b1899 := true;
      b1900 := true;
      b1901 := true;
      b1902 := (b1898 AND (b1899 AND (b1900 AND b1901)));
      b1903 := true;
      r1904 := r1815(0 to 7);
      r1905 := r1815(8 to 15);
      r1906 := r1815(16 to 23);
      r1907 := r1815(24 to 31);
      b1908 := true;
      b1909 := true;
      b1910 := true;
      b1911 := true;
      b1912 := (b1908 AND (b1909 AND (b1910 AND b1911)));
      b1913 := true;
      r1914 := r1816(0 to 7);
      r1915 := r1816(8 to 15);
      r1916 := r1816(16 to 23);
      r1917 := r1816(24 to 31);
      b1918 := true;
      b1919 := true;
      b1920 := true;
      b1921 := true;
      b1922 := (b1918 AND (b1919 AND (b1920 AND b1921)));
      b1923 := true;
      r1924 := r1817(0 to 7);
      r1925 := r1817(8 to 15);
      r1926 := r1817(16 to 23);
      r1927 := r1817(24 to 31);
      b1928 := true;
      b1929 := true;
      b1930 := true;
      b1931 := true;
      b1932 := (b1928 AND (b1929 AND (b1930 AND b1931)));
      b1933 := true;
      r1934 := r1818(0 to 7);
      r1935 := r1818(8 to 15);
      r1936 := r1818(16 to 23);
      r1937 := r1818(24 to 31);
      b1938 := true;
      b1939 := true;
      b1940 := true;
      b1941 := true;
      b1942 := (b1938 AND (b1939 AND (b1940 AND b1941)));
      b1943 := true;
      r1944 := r1819(0 to 7);
      r1945 := r1819(8 to 15);
      r1946 := r1819(16 to 23);
      r1947 := r1819(24 to 31);
      b1948 := true;
      b1949 := true;
      b1950 := true;
      b1951 := true;
      b1952 := (b1948 AND (b1949 AND (b1950 AND b1951)));
      b1953 := true;
      r1954 := r1820(0 to 7);
      r1955 := r1820(8 to 15);
      r1956 := r1820(16 to 23);
      r1957 := r1820(24 to 31);
      b1958 := true;
      b1959 := true;
      b1960 := true;
      b1961 := true;
      b1962 := (b1958 AND (b1959 AND (b1960 AND b1961)));
      b1963 := true;
      r1964 := r1821(0 to 7);
      r1965 := r1821(8 to 15);
      r1966 := r1821(16 to 23);
      r1967 := r1821(24 to 31);
      b1968 := true;
      b1969 := true;
      b1970 := true;
      b1971 := true;
      b1972 := (b1968 AND (b1969 AND (b1970 AND b1971)));
      b1973 := true;
      r1974 := r1822(0 to 7);
      r1975 := r1822(8 to 15);
      r1976 := r1822(16 to 23);
      r1977 := r1822(24 to 31);
      b1978 := true;
      b1979 := true;
      b1980 := true;
      b1981 := true;
      b1982 := (b1978 AND (b1979 AND (b1980 AND b1981)));
      b1983 := (b1832 AND (b1842 AND (b1852 AND (b1862 AND (b1872 AND (b1882 AND (b1892 AND (b1902 AND (b1912 AND (b1922 AND (b1932 AND (b1942 AND (b1952 AND (b1962 AND (b1972 AND b1982)))))))))))))));
      if b1983 then
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        null;
        r1985 := (r1824 & r1825 & r1826 & r1827 & r1834 & r1835 & r1836 & r1837 & r1844 & r1845 & r1846 & r1847 & r1854 & r1855 & r1856 & r1857 & r1864 & r1865 & r1866 & r1867 & r1874 & r1875 & r1876 & r1877 & r1884 & r1885 & r1886 & r1887 & r1894 & r1895 & r1896 & r1897 & r1904 & r1905 & r1906 & r1907 & r1914 & r1915 & r1916 & r1917 & r1924 & r1925 & r1926 & r1927 & r1934 & r1935 & r1936 & r1937 & r1944 & r1945 & r1946 & r1947 & r1954 & r1955 & r1956 & r1957 & r1964 & r1965 & r1966 & r1967 & r1974 & r1975 & r1976 & r1977);
        r1805 := r1985;
      end if;
      r1672 := r1805;
    end if;
    return r1672;
  end rewire_expwords_1669;
  function rewire_littleendianp_1707(r1708 : std_logic_vector) return std_logic_vector
  is
    variable r1786 : std_logic_vector(0 to 31) := (others => '0');
    variable r1785 : std_logic_vector(0 to 7) := (others => '0');
    variable r1783 : std_logic_vector(0 to 7) := (others => '0');
    variable r1781 : std_logic_vector(0 to 7) := (others => '0');
    variable r1779 : std_logic_vector(0 to 7) := (others => '0');
    variable b1776 : boolean := false;
    variable b1775 : boolean := false;
    variable b1774 : boolean := false;
    variable b1773 : boolean := false;
    variable b1772 : boolean := false;
    variable b1771 : boolean := false;
    variable b1770 : boolean := false;
    variable b1769 : boolean := false;
    variable b1768 : boolean := false;
    variable b1767 : boolean := false;
    variable b1766 : boolean := false;
    variable b1765 : boolean := false;
    variable b1764 : boolean := false;
    variable b1763 : boolean := false;
    variable b1762 : boolean := false;
    variable b1761 : boolean := false;
    variable b1760 : boolean := false;
    variable b1759 : boolean := false;
    variable b1758 : boolean := false;
    variable b1757 : boolean := false;
    variable b1756 : boolean := false;
    variable b1755 : boolean := false;
    variable b1754 : boolean := false;
    variable b1753 : boolean := false;
    variable b1752 : boolean := false;
    variable b1751 : boolean := false;
    variable b1750 : boolean := false;
    variable b1749 : boolean := false;
    variable b1748 : boolean := false;
    variable b1747 : boolean := false;
    variable b1746 : boolean := false;
    variable b1745 : boolean := false;
    variable b1744 : boolean := false;
    variable r1743 : std_logic_vector(0 to 0) := (others => '0');
    variable r1742 : std_logic_vector(0 to 0) := (others => '0');
    variable r1741 : std_logic_vector(0 to 0) := (others => '0');
    variable r1740 : std_logic_vector(0 to 0) := (others => '0');
    variable r1739 : std_logic_vector(0 to 0) := (others => '0');
    variable r1738 : std_logic_vector(0 to 0) := (others => '0');
    variable r1737 : std_logic_vector(0 to 0) := (others => '0');
    variable r1736 : std_logic_vector(0 to 0) := (others => '0');
    variable r1735 : std_logic_vector(0 to 0) := (others => '0');
    variable r1734 : std_logic_vector(0 to 0) := (others => '0');
    variable r1733 : std_logic_vector(0 to 0) := (others => '0');
    variable r1732 : std_logic_vector(0 to 0) := (others => '0');
    variable r1731 : std_logic_vector(0 to 0) := (others => '0');
    variable r1730 : std_logic_vector(0 to 0) := (others => '0');
    variable r1729 : std_logic_vector(0 to 0) := (others => '0');
    variable r1728 : std_logic_vector(0 to 0) := (others => '0');
    variable r1727 : std_logic_vector(0 to 0) := (others => '0');
    variable r1726 : std_logic_vector(0 to 0) := (others => '0');
    variable r1725 : std_logic_vector(0 to 0) := (others => '0');
    variable r1724 : std_logic_vector(0 to 0) := (others => '0');
    variable r1723 : std_logic_vector(0 to 0) := (others => '0');
    variable r1722 : std_logic_vector(0 to 0) := (others => '0');
    variable r1721 : std_logic_vector(0 to 0) := (others => '0');
    variable r1720 : std_logic_vector(0 to 0) := (others => '0');
    variable r1719 : std_logic_vector(0 to 0) := (others => '0');
    variable r1718 : std_logic_vector(0 to 0) := (others => '0');
    variable r1717 : std_logic_vector(0 to 0) := (others => '0');
    variable r1716 : std_logic_vector(0 to 0) := (others => '0');
    variable r1715 : std_logic_vector(0 to 0) := (others => '0');
    variable r1714 : std_logic_vector(0 to 0) := (others => '0');
    variable r1713 : std_logic_vector(0 to 0) := (others => '0');
    variable r1712 : std_logic_vector(0 to 0) := (others => '0');
    variable b1711 : boolean := false;
    variable r1710 : std_logic_vector(0 to 31) := (others => '0');
  begin
    b1711 := true;
    r1712 := r1708(0 to 0);
    r1713 := r1708(1 to 1);
    r1714 := r1708(2 to 2);
    r1715 := r1708(3 to 3);
    r1716 := r1708(4 to 4);
    r1717 := r1708(5 to 5);
    r1718 := r1708(6 to 6);
    r1719 := r1708(7 to 7);
    r1720 := r1708(8 to 8);
    r1721 := r1708(9 to 9);
    r1722 := r1708(10 to 10);
    r1723 := r1708(11 to 11);
    r1724 := r1708(12 to 12);
    r1725 := r1708(13 to 13);
    r1726 := r1708(14 to 14);
    r1727 := r1708(15 to 15);
    r1728 := r1708(16 to 16);
    r1729 := r1708(17 to 17);
    r1730 := r1708(18 to 18);
    r1731 := r1708(19 to 19);
    r1732 := r1708(20 to 20);
    r1733 := r1708(21 to 21);
    r1734 := r1708(22 to 22);
    r1735 := r1708(23 to 23);
    r1736 := r1708(24 to 24);
    r1737 := r1708(25 to 25);
    r1738 := r1708(26 to 26);
    r1739 := r1708(27 to 27);
    r1740 := r1708(28 to 28);
    r1741 := r1708(29 to 29);
    r1742 := r1708(30 to 30);
    r1743 := r1708(31 to 31);
    b1744 := true;
    b1745 := true;
    b1746 := true;
    b1747 := true;
    b1748 := true;
    b1749 := true;
    b1750 := true;
    b1751 := true;
    b1752 := true;
    b1753 := true;
    b1754 := true;
    b1755 := true;
    b1756 := true;
    b1757 := true;
    b1758 := true;
    b1759 := true;
    b1760 := true;
    b1761 := true;
    b1762 := true;
    b1763 := true;
    b1764 := true;
    b1765 := true;
    b1766 := true;
    b1767 := true;
    b1768 := true;
    b1769 := true;
    b1770 := true;
    b1771 := true;
    b1772 := true;
    b1773 := true;
    b1774 := true;
    b1775 := true;
    b1776 := (b1744 AND (b1745 AND (b1746 AND (b1747 AND (b1748 AND (b1749 AND (b1750 AND (b1751 AND (b1752 AND (b1753 AND (b1754 AND (b1755 AND (b1756 AND (b1757 AND (b1758 AND (b1759 AND (b1760 AND (b1761 AND (b1762 AND (b1763 AND (b1764 AND (b1765 AND (b1766 AND (b1767 AND (b1768 AND (b1769 AND (b1770 AND (b1771 AND (b1772 AND (b1773 AND (b1774 AND b1775)))))))))))))))))))))))))))))));
    if b1776 then
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      r1779 := (r1736 & r1737 & r1738 & r1739 & r1740 & r1741 & r1742 & r1743);
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      r1781 := (r1728 & r1729 & r1730 & r1731 & r1732 & r1733 & r1734 & r1735);
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      r1783 := (r1720 & r1721 & r1722 & r1723 & r1724 & r1725 & r1726 & r1727);
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      null;
      r1785 := (r1712 & r1713 & r1714 & r1715 & r1716 & r1717 & r1718 & r1719);
      r1786 := (r1779 & r1781 & r1783 & r1785);
      r1710 := r1786;
    end if;
    return r1710;
  end rewire_littleendianp_1707;
  function rewire_sigma3_1541 return std_logic_vector
  is
    variable r1616 : std_logic_vector(0 to 31) := (others => '0');
    variable r1615 : std_logic_vector(0 to 7) := (others => '0');
    variable r1613 : std_logic_vector(0 to 0) := (others => '0');
    variable r1611 : std_logic_vector(0 to 0) := (others => '0');
    variable r1609 : std_logic_vector(0 to 0) := (others => '0');
    variable r1607 : std_logic_vector(0 to 0) := (others => '0');
    variable r1605 : std_logic_vector(0 to 0) := (others => '0');
    variable r1603 : std_logic_vector(0 to 0) := (others => '0');
    variable r1601 : std_logic_vector(0 to 0) := (others => '0');
    variable r1599 : std_logic_vector(0 to 0) := (others => '0');
    variable r1597 : std_logic_vector(0 to 7) := (others => '0');
    variable r1595 : std_logic_vector(0 to 0) := (others => '0');
    variable r1593 : std_logic_vector(0 to 0) := (others => '0');
    variable r1591 : std_logic_vector(0 to 0) := (others => '0');
    variable r1589 : std_logic_vector(0 to 0) := (others => '0');
    variable r1587 : std_logic_vector(0 to 0) := (others => '0');
    variable r1585 : std_logic_vector(0 to 0) := (others => '0');
    variable r1583 : std_logic_vector(0 to 0) := (others => '0');
    variable r1581 : std_logic_vector(0 to 0) := (others => '0');
    variable r1579 : std_logic_vector(0 to 7) := (others => '0');
    variable r1577 : std_logic_vector(0 to 0) := (others => '0');
    variable r1575 : std_logic_vector(0 to 0) := (others => '0');
    variable r1573 : std_logic_vector(0 to 0) := (others => '0');
    variable r1571 : std_logic_vector(0 to 0) := (others => '0');
    variable r1569 : std_logic_vector(0 to 0) := (others => '0');
    variable r1567 : std_logic_vector(0 to 0) := (others => '0');
    variable r1565 : std_logic_vector(0 to 0) := (others => '0');
    variable r1563 : std_logic_vector(0 to 0) := (others => '0');
    variable r1561 : std_logic_vector(0 to 7) := (others => '0');
    variable r1559 : std_logic_vector(0 to 0) := (others => '0');
    variable r1557 : std_logic_vector(0 to 0) := (others => '0');
    variable r1555 : std_logic_vector(0 to 0) := (others => '0');
    variable r1553 : std_logic_vector(0 to 0) := (others => '0');
    variable r1551 : std_logic_vector(0 to 0) := (others => '0');
    variable r1549 : std_logic_vector(0 to 0) := (others => '0');
    variable r1547 : std_logic_vector(0 to 0) := (others => '0');
    variable r1545 : std_logic_vector(0 to 0) := (others => '0');
  begin
    r1545 := "1";
    r1547 := "1";
    r1549 := "0";
    r1551 := "1";
    r1553 := "0";
    r1555 := "0";
    r1557 := "0";
    r1559 := "1";
    r1561 := (r1545 & r1547 & r1549 & r1551 & r1553 & r1555 & r1557 & r1559);
    r1563 := "0";
    r1565 := "1";
    r1567 := "0";
    r1569 := "1";
    r1571 := "1";
    r1573 := "0";
    r1575 := "0";
    r1577 := "1";
    r1579 := (r1563 & r1565 & r1567 & r1569 & r1571 & r1573 & r1575 & r1577);
    r1581 := "1";
    r1583 := "1";
    r1585 := "1";
    r1587 := "1";
    r1589 := "1";
    r1591 := "0";
    r1593 := "1";
    r1595 := "1";
    r1597 := (r1581 & r1583 & r1585 & r1587 & r1589 & r1591 & r1593 & r1595);
    r1599 := "0";
    r1601 := "0";
    r1603 := "1";
    r1605 := "0";
    r1607 := "1";
    r1609 := "0";
    r1611 := "0";
    r1613 := "1";
    r1615 := (r1599 & r1601 & r1603 & r1605 & r1607 & r1609 & r1611 & r1613);
    r1616 := (r1561 & r1579 & r1597 & r1615);
    return r1616;
  end rewire_sigma3_1541;
  function rewire_sigma2_1464 return std_logic_vector
  is
    variable r1539 : std_logic_vector(0 to 31) := (others => '0');
    variable r1538 : std_logic_vector(0 to 7) := (others => '0');
    variable r1536 : std_logic_vector(0 to 0) := (others => '0');
    variable r1534 : std_logic_vector(0 to 0) := (others => '0');
    variable r1532 : std_logic_vector(0 to 0) := (others => '0');
    variable r1530 : std_logic_vector(0 to 0) := (others => '0');
    variable r1528 : std_logic_vector(0 to 0) := (others => '0');
    variable r1526 : std_logic_vector(0 to 0) := (others => '0');
    variable r1524 : std_logic_vector(0 to 0) := (others => '0');
    variable r1522 : std_logic_vector(0 to 0) := (others => '0');
    variable r1520 : std_logic_vector(0 to 7) := (others => '0');
    variable r1518 : std_logic_vector(0 to 0) := (others => '0');
    variable r1516 : std_logic_vector(0 to 0) := (others => '0');
    variable r1514 : std_logic_vector(0 to 0) := (others => '0');
    variable r1512 : std_logic_vector(0 to 0) := (others => '0');
    variable r1510 : std_logic_vector(0 to 0) := (others => '0');
    variable r1508 : std_logic_vector(0 to 0) := (others => '0');
    variable r1506 : std_logic_vector(0 to 0) := (others => '0');
    variable r1504 : std_logic_vector(0 to 0) := (others => '0');
    variable r1502 : std_logic_vector(0 to 7) := (others => '0');
    variable r1500 : std_logic_vector(0 to 0) := (others => '0');
    variable r1498 : std_logic_vector(0 to 0) := (others => '0');
    variable r1496 : std_logic_vector(0 to 0) := (others => '0');
    variable r1494 : std_logic_vector(0 to 0) := (others => '0');
    variable r1492 : std_logic_vector(0 to 0) := (others => '0');
    variable r1490 : std_logic_vector(0 to 0) := (others => '0');
    variable r1488 : std_logic_vector(0 to 0) := (others => '0');
    variable r1486 : std_logic_vector(0 to 0) := (others => '0');
    variable r1484 : std_logic_vector(0 to 7) := (others => '0');
    variable r1482 : std_logic_vector(0 to 0) := (others => '0');
    variable r1480 : std_logic_vector(0 to 0) := (others => '0');
    variable r1478 : std_logic_vector(0 to 0) := (others => '0');
    variable r1476 : std_logic_vector(0 to 0) := (others => '0');
    variable r1474 : std_logic_vector(0 to 0) := (others => '0');
    variable r1472 : std_logic_vector(0 to 0) := (others => '0');
    variable r1470 : std_logic_vector(0 to 0) := (others => '0');
    variable r1468 : std_logic_vector(0 to 0) := (others => '0');
  begin
    r1468 := "1";
    r1470 := "0";
    r1472 := "1";
    r1474 := "1";
    r1476 := "0";
    r1478 := "0";
    r1480 := "1";
    r1482 := "1";
    r1484 := (r1468 & r1470 & r1472 & r1474 & r1476 & r1478 & r1480 & r1482);
    r1486 := "0";
    r1488 := "1";
    r1490 := "0";
    r1492 := "0";
    r1494 := "1";
    r1496 := "0";
    r1498 := "1";
    r1500 := "1";
    r1502 := (r1486 & r1488 & r1490 & r1492 & r1494 & r1496 & r1498 & r1500);
    r1504 := "1";
    r1506 := "0";
    r1508 := "1";
    r1510 := "1";
    r1512 := "1";
    r1514 := "0";
    r1516 := "0";
    r1518 := "1";
    r1520 := (r1504 & r1506 & r1508 & r1510 & r1512 & r1514 & r1516 & r1518);
    r1522 := "0";
    r1524 := "1";
    r1526 := "1";
    r1528 := "0";
    r1530 := "0";
    r1532 := "0";
    r1534 := "0";
    r1536 := "1";
    r1538 := (r1522 & r1524 & r1526 & r1528 & r1530 & r1532 & r1534 & r1536);
    r1539 := (r1484 & r1502 & r1520 & r1538);
    return r1539;
  end rewire_sigma2_1464;
  function rewire_sigma1_1387 return std_logic_vector
  is
    variable r1462 : std_logic_vector(0 to 31) := (others => '0');
    variable r1461 : std_logic_vector(0 to 7) := (others => '0');
    variable r1459 : std_logic_vector(0 to 0) := (others => '0');
    variable r1457 : std_logic_vector(0 to 0) := (others => '0');
    variable r1455 : std_logic_vector(0 to 0) := (others => '0');
    variable r1453 : std_logic_vector(0 to 0) := (others => '0');
    variable r1451 : std_logic_vector(0 to 0) := (others => '0');
    variable r1449 : std_logic_vector(0 to 0) := (others => '0');
    variable r1447 : std_logic_vector(0 to 0) := (others => '0');
    variable r1445 : std_logic_vector(0 to 0) := (others => '0');
    variable r1443 : std_logic_vector(0 to 7) := (others => '0');
    variable r1441 : std_logic_vector(0 to 0) := (others => '0');
    variable r1439 : std_logic_vector(0 to 0) := (others => '0');
    variable r1437 : std_logic_vector(0 to 0) := (others => '0');
    variable r1435 : std_logic_vector(0 to 0) := (others => '0');
    variable r1433 : std_logic_vector(0 to 0) := (others => '0');
    variable r1431 : std_logic_vector(0 to 0) := (others => '0');
    variable r1429 : std_logic_vector(0 to 0) := (others => '0');
    variable r1427 : std_logic_vector(0 to 0) := (others => '0');
    variable r1425 : std_logic_vector(0 to 7) := (others => '0');
    variable r1423 : std_logic_vector(0 to 0) := (others => '0');
    variable r1421 : std_logic_vector(0 to 0) := (others => '0');
    variable r1419 : std_logic_vector(0 to 0) := (others => '0');
    variable r1417 : std_logic_vector(0 to 0) := (others => '0');
    variable r1415 : std_logic_vector(0 to 0) := (others => '0');
    variable r1413 : std_logic_vector(0 to 0) := (others => '0');
    variable r1411 : std_logic_vector(0 to 0) := (others => '0');
    variable r1409 : std_logic_vector(0 to 0) := (others => '0');
    variable r1407 : std_logic_vector(0 to 7) := (others => '0');
    variable r1405 : std_logic_vector(0 to 0) := (others => '0');
    variable r1403 : std_logic_vector(0 to 0) := (others => '0');
    variable r1401 : std_logic_vector(0 to 0) := (others => '0');
    variable r1399 : std_logic_vector(0 to 0) := (others => '0');
    variable r1397 : std_logic_vector(0 to 0) := (others => '0');
    variable r1395 : std_logic_vector(0 to 0) := (others => '0');
    variable r1393 : std_logic_vector(0 to 0) := (others => '0');
    variable r1391 : std_logic_vector(0 to 0) := (others => '0');
  begin
    r1391 := "1";
    r1393 := "0";
    r1395 := "0";
    r1397 := "0";
    r1399 := "1";
    r1401 := "0";
    r1403 := "0";
    r1405 := "1";
    r1407 := (r1391 & r1393 & r1395 & r1397 & r1399 & r1401 & r1403 & r1405);
    r1409 := "1";
    r1411 := "1";
    r1413 := "0";
    r1415 := "1";
    r1417 := "1";
    r1419 := "0";
    r1421 := "0";
    r1423 := "1";
    r1425 := (r1409 & r1411 & r1413 & r1415 & r1417 & r1419 & r1421 & r1423);
    r1427 := "1";
    r1429 := "1";
    r1431 := "1";
    r1433 := "1";
    r1435 := "1";
    r1437 := "0";
    r1439 := "1";
    r1441 := "1";
    r1443 := (r1427 & r1429 & r1431 & r1433 & r1435 & r1437 & r1439 & r1441);
    r1445 := "0";
    r1447 := "0";
    r1449 := "1";
    r1451 := "1";
    r1453 := "0";
    r1455 := "0";
    r1457 := "1";
    r1459 := "1";
    r1461 := (r1445 & r1447 & r1449 & r1451 & r1453 & r1455 & r1457 & r1459);
    r1462 := (r1407 & r1425 & r1443 & r1461);
    return r1462;
  end rewire_sigma1_1387;
  function rewire_sigma0_1310 return std_logic_vector
  is
    variable r1385 : std_logic_vector(0 to 31) := (others => '0');
    variable r1384 : std_logic_vector(0 to 7) := (others => '0');
    variable r1382 : std_logic_vector(0 to 0) := (others => '0');
    variable r1380 : std_logic_vector(0 to 0) := (others => '0');
    variable r1378 : std_logic_vector(0 to 0) := (others => '0');
    variable r1376 : std_logic_vector(0 to 0) := (others => '0');
    variable r1374 : std_logic_vector(0 to 0) := (others => '0');
    variable r1372 : std_logic_vector(0 to 0) := (others => '0');
    variable r1370 : std_logic_vector(0 to 0) := (others => '0');
    variable r1368 : std_logic_vector(0 to 0) := (others => '0');
    variable r1366 : std_logic_vector(0 to 7) := (others => '0');
    variable r1364 : std_logic_vector(0 to 0) := (others => '0');
    variable r1362 : std_logic_vector(0 to 0) := (others => '0');
    variable r1360 : std_logic_vector(0 to 0) := (others => '0');
    variable r1358 : std_logic_vector(0 to 0) := (others => '0');
    variable r1356 : std_logic_vector(0 to 0) := (others => '0');
    variable r1354 : std_logic_vector(0 to 0) := (others => '0');
    variable r1352 : std_logic_vector(0 to 0) := (others => '0');
    variable r1350 : std_logic_vector(0 to 0) := (others => '0');
    variable r1348 : std_logic_vector(0 to 7) := (others => '0');
    variable r1346 : std_logic_vector(0 to 0) := (others => '0');
    variable r1344 : std_logic_vector(0 to 0) := (others => '0');
    variable r1342 : std_logic_vector(0 to 0) := (others => '0');
    variable r1340 : std_logic_vector(0 to 0) := (others => '0');
    variable r1338 : std_logic_vector(0 to 0) := (others => '0');
    variable r1336 : std_logic_vector(0 to 0) := (others => '0');
    variable r1334 : std_logic_vector(0 to 0) := (others => '0');
    variable r1332 : std_logic_vector(0 to 0) := (others => '0');
    variable r1330 : std_logic_vector(0 to 7) := (others => '0');
    variable r1328 : std_logic_vector(0 to 0) := (others => '0');
    variable r1326 : std_logic_vector(0 to 0) := (others => '0');
    variable r1324 : std_logic_vector(0 to 0) := (others => '0');
    variable r1322 : std_logic_vector(0 to 0) := (others => '0');
    variable r1320 : std_logic_vector(0 to 0) := (others => '0');
    variable r1318 : std_logic_vector(0 to 0) := (others => '0');
    variable r1316 : std_logic_vector(0 to 0) := (others => '0');
    variable r1314 : std_logic_vector(0 to 0) := (others => '0');
  begin
    r1314 := "0";
    r1316 := "1";
    r1318 := "0";
    r1320 := "1";
    r1322 := "1";
    r1324 := "0";
    r1326 := "0";
    r1328 := "1";
    r1330 := (r1314 & r1316 & r1318 & r1320 & r1322 & r1324 & r1326 & r1328);
    r1332 := "1";
    r1334 := "1";
    r1336 := "1";
    r1338 := "0";
    r1340 := "0";
    r1342 := "0";
    r1344 := "0";
    r1346 := "1";
    r1348 := (r1332 & r1334 & r1336 & r1338 & r1340 & r1342 & r1344 & r1346);
    r1350 := "1";
    r1352 := "1";
    r1354 := "1";
    r1356 := "1";
    r1358 := "0";
    r1360 := "0";
    r1362 := "0";
    r1364 := "1";
    r1366 := (r1350 & r1352 & r1354 & r1356 & r1358 & r1360 & r1362 & r1364);
    r1368 := "0";
    r1370 := "1";
    r1372 := "1";
    r1374 := "1";
    r1376 := "1";
    r1378 := "0";
    r1380 := "0";
    r1382 := "1";
    r1384 := (r1368 & r1370 & r1372 & r1374 & r1376 & r1378 & r1380 & r1382);
    r1385 := (r1330 & r1348 & r1366 & r1384);
    return r1385;
  end rewire_sigma0_1310;
  function rewire_zerothoutput_3 return std_logic_vector
  is
    variable r1158 : std_logic_vector(0 to 511) := (others => '0');
    variable r1157 : std_logic_vector(0 to 7) := (others => '0');
    variable r1155 : std_logic_vector(0 to 0) := (others => '0');
    variable r1153 : std_logic_vector(0 to 0) := (others => '0');
    variable r1151 : std_logic_vector(0 to 0) := (others => '0');
    variable r1149 : std_logic_vector(0 to 0) := (others => '0');
    variable r1147 : std_logic_vector(0 to 0) := (others => '0');
    variable r1145 : std_logic_vector(0 to 0) := (others => '0');
    variable r1143 : std_logic_vector(0 to 0) := (others => '0');
    variable r1141 : std_logic_vector(0 to 0) := (others => '0');
    variable r1139 : std_logic_vector(0 to 7) := (others => '0');
    variable r1137 : std_logic_vector(0 to 0) := (others => '0');
    variable r1135 : std_logic_vector(0 to 0) := (others => '0');
    variable r1133 : std_logic_vector(0 to 0) := (others => '0');
    variable r1131 : std_logic_vector(0 to 0) := (others => '0');
    variable r1129 : std_logic_vector(0 to 0) := (others => '0');
    variable r1127 : std_logic_vector(0 to 0) := (others => '0');
    variable r1125 : std_logic_vector(0 to 0) := (others => '0');
    variable r1123 : std_logic_vector(0 to 0) := (others => '0');
    variable r1121 : std_logic_vector(0 to 7) := (others => '0');
    variable r1119 : std_logic_vector(0 to 0) := (others => '0');
    variable r1117 : std_logic_vector(0 to 0) := (others => '0');
    variable r1115 : std_logic_vector(0 to 0) := (others => '0');
    variable r1113 : std_logic_vector(0 to 0) := (others => '0');
    variable r1111 : std_logic_vector(0 to 0) := (others => '0');
    variable r1109 : std_logic_vector(0 to 0) := (others => '0');
    variable r1107 : std_logic_vector(0 to 0) := (others => '0');
    variable r1105 : std_logic_vector(0 to 0) := (others => '0');
    variable r1103 : std_logic_vector(0 to 7) := (others => '0');
    variable r1101 : std_logic_vector(0 to 0) := (others => '0');
    variable r1099 : std_logic_vector(0 to 0) := (others => '0');
    variable r1097 : std_logic_vector(0 to 0) := (others => '0');
    variable r1095 : std_logic_vector(0 to 0) := (others => '0');
    variable r1093 : std_logic_vector(0 to 0) := (others => '0');
    variable r1091 : std_logic_vector(0 to 0) := (others => '0');
    variable r1089 : std_logic_vector(0 to 0) := (others => '0');
    variable r1087 : std_logic_vector(0 to 0) := (others => '0');
    variable r1085 : std_logic_vector(0 to 7) := (others => '0');
    variable r1083 : std_logic_vector(0 to 0) := (others => '0');
    variable r1081 : std_logic_vector(0 to 0) := (others => '0');
    variable r1079 : std_logic_vector(0 to 0) := (others => '0');
    variable r1077 : std_logic_vector(0 to 0) := (others => '0');
    variable r1075 : std_logic_vector(0 to 0) := (others => '0');
    variable r1073 : std_logic_vector(0 to 0) := (others => '0');
    variable r1071 : std_logic_vector(0 to 0) := (others => '0');
    variable r1069 : std_logic_vector(0 to 0) := (others => '0');
    variable r1067 : std_logic_vector(0 to 7) := (others => '0');
    variable r1065 : std_logic_vector(0 to 0) := (others => '0');
    variable r1063 : std_logic_vector(0 to 0) := (others => '0');
    variable r1061 : std_logic_vector(0 to 0) := (others => '0');
    variable r1059 : std_logic_vector(0 to 0) := (others => '0');
    variable r1057 : std_logic_vector(0 to 0) := (others => '0');
    variable r1055 : std_logic_vector(0 to 0) := (others => '0');
    variable r1053 : std_logic_vector(0 to 0) := (others => '0');
    variable r1051 : std_logic_vector(0 to 0) := (others => '0');
    variable r1049 : std_logic_vector(0 to 7) := (others => '0');
    variable r1047 : std_logic_vector(0 to 0) := (others => '0');
    variable r1045 : std_logic_vector(0 to 0) := (others => '0');
    variable r1043 : std_logic_vector(0 to 0) := (others => '0');
    variable r1041 : std_logic_vector(0 to 0) := (others => '0');
    variable r1039 : std_logic_vector(0 to 0) := (others => '0');
    variable r1037 : std_logic_vector(0 to 0) := (others => '0');
    variable r1035 : std_logic_vector(0 to 0) := (others => '0');
    variable r1033 : std_logic_vector(0 to 0) := (others => '0');
    variable r1031 : std_logic_vector(0 to 7) := (others => '0');
    variable r1029 : std_logic_vector(0 to 0) := (others => '0');
    variable r1027 : std_logic_vector(0 to 0) := (others => '0');
    variable r1025 : std_logic_vector(0 to 0) := (others => '0');
    variable r1023 : std_logic_vector(0 to 0) := (others => '0');
    variable r1021 : std_logic_vector(0 to 0) := (others => '0');
    variable r1019 : std_logic_vector(0 to 0) := (others => '0');
    variable r1017 : std_logic_vector(0 to 0) := (others => '0');
    variable r1015 : std_logic_vector(0 to 0) := (others => '0');
    variable r1013 : std_logic_vector(0 to 7) := (others => '0');
    variable r1011 : std_logic_vector(0 to 0) := (others => '0');
    variable r1009 : std_logic_vector(0 to 0) := (others => '0');
    variable r1007 : std_logic_vector(0 to 0) := (others => '0');
    variable r1005 : std_logic_vector(0 to 0) := (others => '0');
    variable r1003 : std_logic_vector(0 to 0) := (others => '0');
    variable r1001 : std_logic_vector(0 to 0) := (others => '0');
    variable r999 : std_logic_vector(0 to 0) := (others => '0');
    variable r997 : std_logic_vector(0 to 0) := (others => '0');
    variable r995 : std_logic_vector(0 to 7) := (others => '0');
    variable r993 : std_logic_vector(0 to 0) := (others => '0');
    variable r991 : std_logic_vector(0 to 0) := (others => '0');
    variable r989 : std_logic_vector(0 to 0) := (others => '0');
    variable r987 : std_logic_vector(0 to 0) := (others => '0');
    variable r985 : std_logic_vector(0 to 0) := (others => '0');
    variable r983 : std_logic_vector(0 to 0) := (others => '0');
    variable r981 : std_logic_vector(0 to 0) := (others => '0');
    variable r979 : std_logic_vector(0 to 0) := (others => '0');
    variable r977 : std_logic_vector(0 to 7) := (others => '0');
    variable r975 : std_logic_vector(0 to 0) := (others => '0');
    variable r973 : std_logic_vector(0 to 0) := (others => '0');
    variable r971 : std_logic_vector(0 to 0) := (others => '0');
    variable r969 : std_logic_vector(0 to 0) := (others => '0');
    variable r967 : std_logic_vector(0 to 0) := (others => '0');
    variable r965 : std_logic_vector(0 to 0) := (others => '0');
    variable r963 : std_logic_vector(0 to 0) := (others => '0');
    variable r961 : std_logic_vector(0 to 0) := (others => '0');
    variable r959 : std_logic_vector(0 to 7) := (others => '0');
    variable r957 : std_logic_vector(0 to 0) := (others => '0');
    variable r955 : std_logic_vector(0 to 0) := (others => '0');
    variable r953 : std_logic_vector(0 to 0) := (others => '0');
    variable r951 : std_logic_vector(0 to 0) := (others => '0');
    variable r949 : std_logic_vector(0 to 0) := (others => '0');
    variable r947 : std_logic_vector(0 to 0) := (others => '0');
    variable r945 : std_logic_vector(0 to 0) := (others => '0');
    variable r943 : std_logic_vector(0 to 0) := (others => '0');
    variable r941 : std_logic_vector(0 to 7) := (others => '0');
    variable r939 : std_logic_vector(0 to 0) := (others => '0');
    variable r937 : std_logic_vector(0 to 0) := (others => '0');
    variable r935 : std_logic_vector(0 to 0) := (others => '0');
    variable r933 : std_logic_vector(0 to 0) := (others => '0');
    variable r931 : std_logic_vector(0 to 0) := (others => '0');
    variable r929 : std_logic_vector(0 to 0) := (others => '0');
    variable r927 : std_logic_vector(0 to 0) := (others => '0');
    variable r925 : std_logic_vector(0 to 0) := (others => '0');
    variable r923 : std_logic_vector(0 to 7) := (others => '0');
    variable r921 : std_logic_vector(0 to 0) := (others => '0');
    variable r919 : std_logic_vector(0 to 0) := (others => '0');
    variable r917 : std_logic_vector(0 to 0) := (others => '0');
    variable r915 : std_logic_vector(0 to 0) := (others => '0');
    variable r913 : std_logic_vector(0 to 0) := (others => '0');
    variable r911 : std_logic_vector(0 to 0) := (others => '0');
    variable r909 : std_logic_vector(0 to 0) := (others => '0');
    variable r907 : std_logic_vector(0 to 0) := (others => '0');
    variable r905 : std_logic_vector(0 to 7) := (others => '0');
    variable r903 : std_logic_vector(0 to 0) := (others => '0');
    variable r901 : std_logic_vector(0 to 0) := (others => '0');
    variable r899 : std_logic_vector(0 to 0) := (others => '0');
    variable r897 : std_logic_vector(0 to 0) := (others => '0');
    variable r895 : std_logic_vector(0 to 0) := (others => '0');
    variable r893 : std_logic_vector(0 to 0) := (others => '0');
    variable r891 : std_logic_vector(0 to 0) := (others => '0');
    variable r889 : std_logic_vector(0 to 0) := (others => '0');
    variable r887 : std_logic_vector(0 to 7) := (others => '0');
    variable r885 : std_logic_vector(0 to 0) := (others => '0');
    variable r883 : std_logic_vector(0 to 0) := (others => '0');
    variable r881 : std_logic_vector(0 to 0) := (others => '0');
    variable r879 : std_logic_vector(0 to 0) := (others => '0');
    variable r877 : std_logic_vector(0 to 0) := (others => '0');
    variable r875 : std_logic_vector(0 to 0) := (others => '0');
    variable r873 : std_logic_vector(0 to 0) := (others => '0');
    variable r871 : std_logic_vector(0 to 0) := (others => '0');
    variable r869 : std_logic_vector(0 to 7) := (others => '0');
    variable r867 : std_logic_vector(0 to 0) := (others => '0');
    variable r865 : std_logic_vector(0 to 0) := (others => '0');
    variable r863 : std_logic_vector(0 to 0) := (others => '0');
    variable r861 : std_logic_vector(0 to 0) := (others => '0');
    variable r859 : std_logic_vector(0 to 0) := (others => '0');
    variable r857 : std_logic_vector(0 to 0) := (others => '0');
    variable r855 : std_logic_vector(0 to 0) := (others => '0');
    variable r853 : std_logic_vector(0 to 0) := (others => '0');
    variable r851 : std_logic_vector(0 to 7) := (others => '0');
    variable r849 : std_logic_vector(0 to 0) := (others => '0');
    variable r847 : std_logic_vector(0 to 0) := (others => '0');
    variable r845 : std_logic_vector(0 to 0) := (others => '0');
    variable r843 : std_logic_vector(0 to 0) := (others => '0');
    variable r841 : std_logic_vector(0 to 0) := (others => '0');
    variable r839 : std_logic_vector(0 to 0) := (others => '0');
    variable r837 : std_logic_vector(0 to 0) := (others => '0');
    variable r835 : std_logic_vector(0 to 0) := (others => '0');
    variable r833 : std_logic_vector(0 to 7) := (others => '0');
    variable r831 : std_logic_vector(0 to 0) := (others => '0');
    variable r829 : std_logic_vector(0 to 0) := (others => '0');
    variable r827 : std_logic_vector(0 to 0) := (others => '0');
    variable r825 : std_logic_vector(0 to 0) := (others => '0');
    variable r823 : std_logic_vector(0 to 0) := (others => '0');
    variable r821 : std_logic_vector(0 to 0) := (others => '0');
    variable r819 : std_logic_vector(0 to 0) := (others => '0');
    variable r817 : std_logic_vector(0 to 0) := (others => '0');
    variable r815 : std_logic_vector(0 to 7) := (others => '0');
    variable r813 : std_logic_vector(0 to 0) := (others => '0');
    variable r811 : std_logic_vector(0 to 0) := (others => '0');
    variable r809 : std_logic_vector(0 to 0) := (others => '0');
    variable r807 : std_logic_vector(0 to 0) := (others => '0');
    variable r805 : std_logic_vector(0 to 0) := (others => '0');
    variable r803 : std_logic_vector(0 to 0) := (others => '0');
    variable r801 : std_logic_vector(0 to 0) := (others => '0');
    variable r799 : std_logic_vector(0 to 0) := (others => '0');
    variable r797 : std_logic_vector(0 to 7) := (others => '0');
    variable r795 : std_logic_vector(0 to 0) := (others => '0');
    variable r793 : std_logic_vector(0 to 0) := (others => '0');
    variable r791 : std_logic_vector(0 to 0) := (others => '0');
    variable r789 : std_logic_vector(0 to 0) := (others => '0');
    variable r787 : std_logic_vector(0 to 0) := (others => '0');
    variable r785 : std_logic_vector(0 to 0) := (others => '0');
    variable r783 : std_logic_vector(0 to 0) := (others => '0');
    variable r781 : std_logic_vector(0 to 0) := (others => '0');
    variable r779 : std_logic_vector(0 to 7) := (others => '0');
    variable r777 : std_logic_vector(0 to 0) := (others => '0');
    variable r775 : std_logic_vector(0 to 0) := (others => '0');
    variable r773 : std_logic_vector(0 to 0) := (others => '0');
    variable r771 : std_logic_vector(0 to 0) := (others => '0');
    variable r769 : std_logic_vector(0 to 0) := (others => '0');
    variable r767 : std_logic_vector(0 to 0) := (others => '0');
    variable r765 : std_logic_vector(0 to 0) := (others => '0');
    variable r763 : std_logic_vector(0 to 0) := (others => '0');
    variable r761 : std_logic_vector(0 to 7) := (others => '0');
    variable r759 : std_logic_vector(0 to 0) := (others => '0');
    variable r757 : std_logic_vector(0 to 0) := (others => '0');
    variable r755 : std_logic_vector(0 to 0) := (others => '0');
    variable r753 : std_logic_vector(0 to 0) := (others => '0');
    variable r751 : std_logic_vector(0 to 0) := (others => '0');
    variable r749 : std_logic_vector(0 to 0) := (others => '0');
    variable r747 : std_logic_vector(0 to 0) := (others => '0');
    variable r745 : std_logic_vector(0 to 0) := (others => '0');
    variable r743 : std_logic_vector(0 to 7) := (others => '0');
    variable r741 : std_logic_vector(0 to 0) := (others => '0');
    variable r739 : std_logic_vector(0 to 0) := (others => '0');
    variable r737 : std_logic_vector(0 to 0) := (others => '0');
    variable r735 : std_logic_vector(0 to 0) := (others => '0');
    variable r733 : std_logic_vector(0 to 0) := (others => '0');
    variable r731 : std_logic_vector(0 to 0) := (others => '0');
    variable r729 : std_logic_vector(0 to 0) := (others => '0');
    variable r727 : std_logic_vector(0 to 0) := (others => '0');
    variable r725 : std_logic_vector(0 to 7) := (others => '0');
    variable r723 : std_logic_vector(0 to 0) := (others => '0');
    variable r721 : std_logic_vector(0 to 0) := (others => '0');
    variable r719 : std_logic_vector(0 to 0) := (others => '0');
    variable r717 : std_logic_vector(0 to 0) := (others => '0');
    variable r715 : std_logic_vector(0 to 0) := (others => '0');
    variable r713 : std_logic_vector(0 to 0) := (others => '0');
    variable r711 : std_logic_vector(0 to 0) := (others => '0');
    variable r709 : std_logic_vector(0 to 0) := (others => '0');
    variable r707 : std_logic_vector(0 to 7) := (others => '0');
    variable r705 : std_logic_vector(0 to 0) := (others => '0');
    variable r703 : std_logic_vector(0 to 0) := (others => '0');
    variable r701 : std_logic_vector(0 to 0) := (others => '0');
    variable r699 : std_logic_vector(0 to 0) := (others => '0');
    variable r697 : std_logic_vector(0 to 0) := (others => '0');
    variable r695 : std_logic_vector(0 to 0) := (others => '0');
    variable r693 : std_logic_vector(0 to 0) := (others => '0');
    variable r691 : std_logic_vector(0 to 0) := (others => '0');
    variable r689 : std_logic_vector(0 to 7) := (others => '0');
    variable r687 : std_logic_vector(0 to 0) := (others => '0');
    variable r685 : std_logic_vector(0 to 0) := (others => '0');
    variable r683 : std_logic_vector(0 to 0) := (others => '0');
    variable r681 : std_logic_vector(0 to 0) := (others => '0');
    variable r679 : std_logic_vector(0 to 0) := (others => '0');
    variable r677 : std_logic_vector(0 to 0) := (others => '0');
    variable r675 : std_logic_vector(0 to 0) := (others => '0');
    variable r673 : std_logic_vector(0 to 0) := (others => '0');
    variable r671 : std_logic_vector(0 to 7) := (others => '0');
    variable r669 : std_logic_vector(0 to 0) := (others => '0');
    variable r667 : std_logic_vector(0 to 0) := (others => '0');
    variable r665 : std_logic_vector(0 to 0) := (others => '0');
    variable r663 : std_logic_vector(0 to 0) := (others => '0');
    variable r661 : std_logic_vector(0 to 0) := (others => '0');
    variable r659 : std_logic_vector(0 to 0) := (others => '0');
    variable r657 : std_logic_vector(0 to 0) := (others => '0');
    variable r655 : std_logic_vector(0 to 0) := (others => '0');
    variable r653 : std_logic_vector(0 to 7) := (others => '0');
    variable r651 : std_logic_vector(0 to 0) := (others => '0');
    variable r649 : std_logic_vector(0 to 0) := (others => '0');
    variable r647 : std_logic_vector(0 to 0) := (others => '0');
    variable r645 : std_logic_vector(0 to 0) := (others => '0');
    variable r643 : std_logic_vector(0 to 0) := (others => '0');
    variable r641 : std_logic_vector(0 to 0) := (others => '0');
    variable r639 : std_logic_vector(0 to 0) := (others => '0');
    variable r637 : std_logic_vector(0 to 0) := (others => '0');
    variable r635 : std_logic_vector(0 to 7) := (others => '0');
    variable r633 : std_logic_vector(0 to 0) := (others => '0');
    variable r631 : std_logic_vector(0 to 0) := (others => '0');
    variable r629 : std_logic_vector(0 to 0) := (others => '0');
    variable r627 : std_logic_vector(0 to 0) := (others => '0');
    variable r625 : std_logic_vector(0 to 0) := (others => '0');
    variable r623 : std_logic_vector(0 to 0) := (others => '0');
    variable r621 : std_logic_vector(0 to 0) := (others => '0');
    variable r619 : std_logic_vector(0 to 0) := (others => '0');
    variable r617 : std_logic_vector(0 to 7) := (others => '0');
    variable r615 : std_logic_vector(0 to 0) := (others => '0');
    variable r613 : std_logic_vector(0 to 0) := (others => '0');
    variable r611 : std_logic_vector(0 to 0) := (others => '0');
    variable r609 : std_logic_vector(0 to 0) := (others => '0');
    variable r607 : std_logic_vector(0 to 0) := (others => '0');
    variable r605 : std_logic_vector(0 to 0) := (others => '0');
    variable r603 : std_logic_vector(0 to 0) := (others => '0');
    variable r601 : std_logic_vector(0 to 0) := (others => '0');
    variable r599 : std_logic_vector(0 to 7) := (others => '0');
    variable r597 : std_logic_vector(0 to 0) := (others => '0');
    variable r595 : std_logic_vector(0 to 0) := (others => '0');
    variable r593 : std_logic_vector(0 to 0) := (others => '0');
    variable r591 : std_logic_vector(0 to 0) := (others => '0');
    variable r589 : std_logic_vector(0 to 0) := (others => '0');
    variable r587 : std_logic_vector(0 to 0) := (others => '0');
    variable r585 : std_logic_vector(0 to 0) := (others => '0');
    variable r583 : std_logic_vector(0 to 0) := (others => '0');
    variable r581 : std_logic_vector(0 to 7) := (others => '0');
    variable r579 : std_logic_vector(0 to 0) := (others => '0');
    variable r577 : std_logic_vector(0 to 0) := (others => '0');
    variable r575 : std_logic_vector(0 to 0) := (others => '0');
    variable r573 : std_logic_vector(0 to 0) := (others => '0');
    variable r571 : std_logic_vector(0 to 0) := (others => '0');
    variable r569 : std_logic_vector(0 to 0) := (others => '0');
    variable r567 : std_logic_vector(0 to 0) := (others => '0');
    variable r565 : std_logic_vector(0 to 0) := (others => '0');
    variable r563 : std_logic_vector(0 to 7) := (others => '0');
    variable r561 : std_logic_vector(0 to 0) := (others => '0');
    variable r559 : std_logic_vector(0 to 0) := (others => '0');
    variable r557 : std_logic_vector(0 to 0) := (others => '0');
    variable r555 : std_logic_vector(0 to 0) := (others => '0');
    variable r553 : std_logic_vector(0 to 0) := (others => '0');
    variable r551 : std_logic_vector(0 to 0) := (others => '0');
    variable r549 : std_logic_vector(0 to 0) := (others => '0');
    variable r547 : std_logic_vector(0 to 0) := (others => '0');
    variable r545 : std_logic_vector(0 to 7) := (others => '0');
    variable r543 : std_logic_vector(0 to 0) := (others => '0');
    variable r541 : std_logic_vector(0 to 0) := (others => '0');
    variable r539 : std_logic_vector(0 to 0) := (others => '0');
    variable r537 : std_logic_vector(0 to 0) := (others => '0');
    variable r535 : std_logic_vector(0 to 0) := (others => '0');
    variable r533 : std_logic_vector(0 to 0) := (others => '0');
    variable r531 : std_logic_vector(0 to 0) := (others => '0');
    variable r529 : std_logic_vector(0 to 0) := (others => '0');
    variable r527 : std_logic_vector(0 to 7) := (others => '0');
    variable r525 : std_logic_vector(0 to 0) := (others => '0');
    variable r523 : std_logic_vector(0 to 0) := (others => '0');
    variable r521 : std_logic_vector(0 to 0) := (others => '0');
    variable r519 : std_logic_vector(0 to 0) := (others => '0');
    variable r517 : std_logic_vector(0 to 0) := (others => '0');
    variable r515 : std_logic_vector(0 to 0) := (others => '0');
    variable r513 : std_logic_vector(0 to 0) := (others => '0');
    variable r511 : std_logic_vector(0 to 0) := (others => '0');
    variable r509 : std_logic_vector(0 to 7) := (others => '0');
    variable r507 : std_logic_vector(0 to 0) := (others => '0');
    variable r505 : std_logic_vector(0 to 0) := (others => '0');
    variable r503 : std_logic_vector(0 to 0) := (others => '0');
    variable r501 : std_logic_vector(0 to 0) := (others => '0');
    variable r499 : std_logic_vector(0 to 0) := (others => '0');
    variable r497 : std_logic_vector(0 to 0) := (others => '0');
    variable r495 : std_logic_vector(0 to 0) := (others => '0');
    variable r493 : std_logic_vector(0 to 0) := (others => '0');
    variable r491 : std_logic_vector(0 to 7) := (others => '0');
    variable r489 : std_logic_vector(0 to 0) := (others => '0');
    variable r487 : std_logic_vector(0 to 0) := (others => '0');
    variable r485 : std_logic_vector(0 to 0) := (others => '0');
    variable r483 : std_logic_vector(0 to 0) := (others => '0');
    variable r481 : std_logic_vector(0 to 0) := (others => '0');
    variable r479 : std_logic_vector(0 to 0) := (others => '0');
    variable r477 : std_logic_vector(0 to 0) := (others => '0');
    variable r475 : std_logic_vector(0 to 0) := (others => '0');
    variable r473 : std_logic_vector(0 to 7) := (others => '0');
    variable r471 : std_logic_vector(0 to 0) := (others => '0');
    variable r469 : std_logic_vector(0 to 0) := (others => '0');
    variable r467 : std_logic_vector(0 to 0) := (others => '0');
    variable r465 : std_logic_vector(0 to 0) := (others => '0');
    variable r463 : std_logic_vector(0 to 0) := (others => '0');
    variable r461 : std_logic_vector(0 to 0) := (others => '0');
    variable r459 : std_logic_vector(0 to 0) := (others => '0');
    variable r457 : std_logic_vector(0 to 0) := (others => '0');
    variable r455 : std_logic_vector(0 to 7) := (others => '0');
    variable r453 : std_logic_vector(0 to 0) := (others => '0');
    variable r451 : std_logic_vector(0 to 0) := (others => '0');
    variable r449 : std_logic_vector(0 to 0) := (others => '0');
    variable r447 : std_logic_vector(0 to 0) := (others => '0');
    variable r445 : std_logic_vector(0 to 0) := (others => '0');
    variable r443 : std_logic_vector(0 to 0) := (others => '0');
    variable r441 : std_logic_vector(0 to 0) := (others => '0');
    variable r439 : std_logic_vector(0 to 0) := (others => '0');
    variable r437 : std_logic_vector(0 to 7) := (others => '0');
    variable r435 : std_logic_vector(0 to 0) := (others => '0');
    variable r433 : std_logic_vector(0 to 0) := (others => '0');
    variable r431 : std_logic_vector(0 to 0) := (others => '0');
    variable r429 : std_logic_vector(0 to 0) := (others => '0');
    variable r427 : std_logic_vector(0 to 0) := (others => '0');
    variable r425 : std_logic_vector(0 to 0) := (others => '0');
    variable r423 : std_logic_vector(0 to 0) := (others => '0');
    variable r421 : std_logic_vector(0 to 0) := (others => '0');
    variable r419 : std_logic_vector(0 to 7) := (others => '0');
    variable r417 : std_logic_vector(0 to 0) := (others => '0');
    variable r415 : std_logic_vector(0 to 0) := (others => '0');
    variable r413 : std_logic_vector(0 to 0) := (others => '0');
    variable r411 : std_logic_vector(0 to 0) := (others => '0');
    variable r409 : std_logic_vector(0 to 0) := (others => '0');
    variable r407 : std_logic_vector(0 to 0) := (others => '0');
    variable r405 : std_logic_vector(0 to 0) := (others => '0');
    variable r403 : std_logic_vector(0 to 0) := (others => '0');
    variable r401 : std_logic_vector(0 to 7) := (others => '0');
    variable r399 : std_logic_vector(0 to 0) := (others => '0');
    variable r397 : std_logic_vector(0 to 0) := (others => '0');
    variable r395 : std_logic_vector(0 to 0) := (others => '0');
    variable r393 : std_logic_vector(0 to 0) := (others => '0');
    variable r391 : std_logic_vector(0 to 0) := (others => '0');
    variable r389 : std_logic_vector(0 to 0) := (others => '0');
    variable r387 : std_logic_vector(0 to 0) := (others => '0');
    variable r385 : std_logic_vector(0 to 0) := (others => '0');
    variable r383 : std_logic_vector(0 to 7) := (others => '0');
    variable r381 : std_logic_vector(0 to 0) := (others => '0');
    variable r379 : std_logic_vector(0 to 0) := (others => '0');
    variable r377 : std_logic_vector(0 to 0) := (others => '0');
    variable r375 : std_logic_vector(0 to 0) := (others => '0');
    variable r373 : std_logic_vector(0 to 0) := (others => '0');
    variable r371 : std_logic_vector(0 to 0) := (others => '0');
    variable r369 : std_logic_vector(0 to 0) := (others => '0');
    variable r367 : std_logic_vector(0 to 0) := (others => '0');
    variable r365 : std_logic_vector(0 to 7) := (others => '0');
    variable r363 : std_logic_vector(0 to 0) := (others => '0');
    variable r361 : std_logic_vector(0 to 0) := (others => '0');
    variable r359 : std_logic_vector(0 to 0) := (others => '0');
    variable r357 : std_logic_vector(0 to 0) := (others => '0');
    variable r355 : std_logic_vector(0 to 0) := (others => '0');
    variable r353 : std_logic_vector(0 to 0) := (others => '0');
    variable r351 : std_logic_vector(0 to 0) := (others => '0');
    variable r349 : std_logic_vector(0 to 0) := (others => '0');
    variable r347 : std_logic_vector(0 to 7) := (others => '0');
    variable r345 : std_logic_vector(0 to 0) := (others => '0');
    variable r343 : std_logic_vector(0 to 0) := (others => '0');
    variable r341 : std_logic_vector(0 to 0) := (others => '0');
    variable r339 : std_logic_vector(0 to 0) := (others => '0');
    variable r337 : std_logic_vector(0 to 0) := (others => '0');
    variable r335 : std_logic_vector(0 to 0) := (others => '0');
    variable r333 : std_logic_vector(0 to 0) := (others => '0');
    variable r331 : std_logic_vector(0 to 0) := (others => '0');
    variable r329 : std_logic_vector(0 to 7) := (others => '0');
    variable r327 : std_logic_vector(0 to 0) := (others => '0');
    variable r325 : std_logic_vector(0 to 0) := (others => '0');
    variable r323 : std_logic_vector(0 to 0) := (others => '0');
    variable r321 : std_logic_vector(0 to 0) := (others => '0');
    variable r319 : std_logic_vector(0 to 0) := (others => '0');
    variable r317 : std_logic_vector(0 to 0) := (others => '0');
    variable r315 : std_logic_vector(0 to 0) := (others => '0');
    variable r313 : std_logic_vector(0 to 0) := (others => '0');
    variable r311 : std_logic_vector(0 to 7) := (others => '0');
    variable r309 : std_logic_vector(0 to 0) := (others => '0');
    variable r307 : std_logic_vector(0 to 0) := (others => '0');
    variable r305 : std_logic_vector(0 to 0) := (others => '0');
    variable r303 : std_logic_vector(0 to 0) := (others => '0');
    variable r301 : std_logic_vector(0 to 0) := (others => '0');
    variable r299 : std_logic_vector(0 to 0) := (others => '0');
    variable r297 : std_logic_vector(0 to 0) := (others => '0');
    variable r295 : std_logic_vector(0 to 0) := (others => '0');
    variable r293 : std_logic_vector(0 to 7) := (others => '0');
    variable r291 : std_logic_vector(0 to 0) := (others => '0');
    variable r289 : std_logic_vector(0 to 0) := (others => '0');
    variable r287 : std_logic_vector(0 to 0) := (others => '0');
    variable r285 : std_logic_vector(0 to 0) := (others => '0');
    variable r283 : std_logic_vector(0 to 0) := (others => '0');
    variable r281 : std_logic_vector(0 to 0) := (others => '0');
    variable r279 : std_logic_vector(0 to 0) := (others => '0');
    variable r277 : std_logic_vector(0 to 0) := (others => '0');
    variable r275 : std_logic_vector(0 to 7) := (others => '0');
    variable r273 : std_logic_vector(0 to 0) := (others => '0');
    variable r271 : std_logic_vector(0 to 0) := (others => '0');
    variable r269 : std_logic_vector(0 to 0) := (others => '0');
    variable r267 : std_logic_vector(0 to 0) := (others => '0');
    variable r265 : std_logic_vector(0 to 0) := (others => '0');
    variable r263 : std_logic_vector(0 to 0) := (others => '0');
    variable r261 : std_logic_vector(0 to 0) := (others => '0');
    variable r259 : std_logic_vector(0 to 0) := (others => '0');
    variable r257 : std_logic_vector(0 to 7) := (others => '0');
    variable r255 : std_logic_vector(0 to 0) := (others => '0');
    variable r253 : std_logic_vector(0 to 0) := (others => '0');
    variable r251 : std_logic_vector(0 to 0) := (others => '0');
    variable r249 : std_logic_vector(0 to 0) := (others => '0');
    variable r247 : std_logic_vector(0 to 0) := (others => '0');
    variable r245 : std_logic_vector(0 to 0) := (others => '0');
    variable r243 : std_logic_vector(0 to 0) := (others => '0');
    variable r241 : std_logic_vector(0 to 0) := (others => '0');
    variable r239 : std_logic_vector(0 to 7) := (others => '0');
    variable r237 : std_logic_vector(0 to 0) := (others => '0');
    variable r235 : std_logic_vector(0 to 0) := (others => '0');
    variable r233 : std_logic_vector(0 to 0) := (others => '0');
    variable r231 : std_logic_vector(0 to 0) := (others => '0');
    variable r229 : std_logic_vector(0 to 0) := (others => '0');
    variable r227 : std_logic_vector(0 to 0) := (others => '0');
    variable r225 : std_logic_vector(0 to 0) := (others => '0');
    variable r223 : std_logic_vector(0 to 0) := (others => '0');
    variable r221 : std_logic_vector(0 to 7) := (others => '0');
    variable r219 : std_logic_vector(0 to 0) := (others => '0');
    variable r217 : std_logic_vector(0 to 0) := (others => '0');
    variable r215 : std_logic_vector(0 to 0) := (others => '0');
    variable r213 : std_logic_vector(0 to 0) := (others => '0');
    variable r211 : std_logic_vector(0 to 0) := (others => '0');
    variable r209 : std_logic_vector(0 to 0) := (others => '0');
    variable r207 : std_logic_vector(0 to 0) := (others => '0');
    variable r205 : std_logic_vector(0 to 0) := (others => '0');
    variable r203 : std_logic_vector(0 to 7) := (others => '0');
    variable r201 : std_logic_vector(0 to 0) := (others => '0');
    variable r199 : std_logic_vector(0 to 0) := (others => '0');
    variable r197 : std_logic_vector(0 to 0) := (others => '0');
    variable r195 : std_logic_vector(0 to 0) := (others => '0');
    variable r193 : std_logic_vector(0 to 0) := (others => '0');
    variable r191 : std_logic_vector(0 to 0) := (others => '0');
    variable r189 : std_logic_vector(0 to 0) := (others => '0');
    variable r187 : std_logic_vector(0 to 0) := (others => '0');
    variable r185 : std_logic_vector(0 to 7) := (others => '0');
    variable r183 : std_logic_vector(0 to 0) := (others => '0');
    variable r181 : std_logic_vector(0 to 0) := (others => '0');
    variable r179 : std_logic_vector(0 to 0) := (others => '0');
    variable r177 : std_logic_vector(0 to 0) := (others => '0');
    variable r175 : std_logic_vector(0 to 0) := (others => '0');
    variable r173 : std_logic_vector(0 to 0) := (others => '0');
    variable r171 : std_logic_vector(0 to 0) := (others => '0');
    variable r169 : std_logic_vector(0 to 0) := (others => '0');
    variable r167 : std_logic_vector(0 to 7) := (others => '0');
    variable r165 : std_logic_vector(0 to 0) := (others => '0');
    variable r163 : std_logic_vector(0 to 0) := (others => '0');
    variable r161 : std_logic_vector(0 to 0) := (others => '0');
    variable r159 : std_logic_vector(0 to 0) := (others => '0');
    variable r157 : std_logic_vector(0 to 0) := (others => '0');
    variable r155 : std_logic_vector(0 to 0) := (others => '0');
    variable r153 : std_logic_vector(0 to 0) := (others => '0');
    variable r151 : std_logic_vector(0 to 0) := (others => '0');
    variable r149 : std_logic_vector(0 to 7) := (others => '0');
    variable r147 : std_logic_vector(0 to 0) := (others => '0');
    variable r145 : std_logic_vector(0 to 0) := (others => '0');
    variable r143 : std_logic_vector(0 to 0) := (others => '0');
    variable r141 : std_logic_vector(0 to 0) := (others => '0');
    variable r139 : std_logic_vector(0 to 0) := (others => '0');
    variable r137 : std_logic_vector(0 to 0) := (others => '0');
    variable r135 : std_logic_vector(0 to 0) := (others => '0');
    variable r133 : std_logic_vector(0 to 0) := (others => '0');
    variable r131 : std_logic_vector(0 to 7) := (others => '0');
    variable r129 : std_logic_vector(0 to 0) := (others => '0');
    variable r127 : std_logic_vector(0 to 0) := (others => '0');
    variable r125 : std_logic_vector(0 to 0) := (others => '0');
    variable r123 : std_logic_vector(0 to 0) := (others => '0');
    variable r121 : std_logic_vector(0 to 0) := (others => '0');
    variable r119 : std_logic_vector(0 to 0) := (others => '0');
    variable r117 : std_logic_vector(0 to 0) := (others => '0');
    variable r115 : std_logic_vector(0 to 0) := (others => '0');
    variable r113 : std_logic_vector(0 to 7) := (others => '0');
    variable r111 : std_logic_vector(0 to 0) := (others => '0');
    variable r109 : std_logic_vector(0 to 0) := (others => '0');
    variable r107 : std_logic_vector(0 to 0) := (others => '0');
    variable r105 : std_logic_vector(0 to 0) := (others => '0');
    variable r103 : std_logic_vector(0 to 0) := (others => '0');
    variable r101 : std_logic_vector(0 to 0) := (others => '0');
    variable r99 : std_logic_vector(0 to 0) := (others => '0');
    variable r97 : std_logic_vector(0 to 0) := (others => '0');
    variable r95 : std_logic_vector(0 to 7) := (others => '0');
    variable r93 : std_logic_vector(0 to 0) := (others => '0');
    variable r91 : std_logic_vector(0 to 0) := (others => '0');
    variable r89 : std_logic_vector(0 to 0) := (others => '0');
    variable r87 : std_logic_vector(0 to 0) := (others => '0');
    variable r85 : std_logic_vector(0 to 0) := (others => '0');
    variable r83 : std_logic_vector(0 to 0) := (others => '0');
    variable r81 : std_logic_vector(0 to 0) := (others => '0');
    variable r79 : std_logic_vector(0 to 0) := (others => '0');
    variable r77 : std_logic_vector(0 to 7) := (others => '0');
    variable r75 : std_logic_vector(0 to 0) := (others => '0');
    variable r73 : std_logic_vector(0 to 0) := (others => '0');
    variable r71 : std_logic_vector(0 to 0) := (others => '0');
    variable r69 : std_logic_vector(0 to 0) := (others => '0');
    variable r67 : std_logic_vector(0 to 0) := (others => '0');
    variable r65 : std_logic_vector(0 to 0) := (others => '0');
    variable r63 : std_logic_vector(0 to 0) := (others => '0');
    variable r61 : std_logic_vector(0 to 0) := (others => '0');
    variable r59 : std_logic_vector(0 to 7) := (others => '0');
    variable r57 : std_logic_vector(0 to 0) := (others => '0');
    variable r55 : std_logic_vector(0 to 0) := (others => '0');
    variable r53 : std_logic_vector(0 to 0) := (others => '0');
    variable r51 : std_logic_vector(0 to 0) := (others => '0');
    variable r49 : std_logic_vector(0 to 0) := (others => '0');
    variable r47 : std_logic_vector(0 to 0) := (others => '0');
    variable r45 : std_logic_vector(0 to 0) := (others => '0');
    variable r43 : std_logic_vector(0 to 0) := (others => '0');
    variable r41 : std_logic_vector(0 to 7) := (others => '0');
    variable r39 : std_logic_vector(0 to 0) := (others => '0');
    variable r37 : std_logic_vector(0 to 0) := (others => '0');
    variable r35 : std_logic_vector(0 to 0) := (others => '0');
    variable r33 : std_logic_vector(0 to 0) := (others => '0');
    variable r31 : std_logic_vector(0 to 0) := (others => '0');
    variable r29 : std_logic_vector(0 to 0) := (others => '0');
    variable r27 : std_logic_vector(0 to 0) := (others => '0');
    variable r25 : std_logic_vector(0 to 0) := (others => '0');
    variable r23 : std_logic_vector(0 to 7) := (others => '0');
    variable r21 : std_logic_vector(0 to 0) := (others => '0');
    variable r19 : std_logic_vector(0 to 0) := (others => '0');
    variable r17 : std_logic_vector(0 to 0) := (others => '0');
    variable r15 : std_logic_vector(0 to 0) := (others => '0');
    variable r13 : std_logic_vector(0 to 0) := (others => '0');
    variable r11 : std_logic_vector(0 to 0) := (others => '0');
    variable r9 : std_logic_vector(0 to 0) := (others => '0');
    variable r7 : std_logic_vector(0 to 0) := (others => '0');
  begin
    r7 := "1";
    r9 := "1";
    r11 := "1";
    r13 := "1";
    r15 := "1";
    r17 := "1";
    r19 := "1";
    r21 := "1";
    r23 := (r7 & r9 & r11 & r13 & r15 & r17 & r19 & r21);
    r25 := "1";
    r27 := "1";
    r29 := "1";
    r31 := "1";
    r33 := "1";
    r35 := "1";
    r37 := "1";
    r39 := "1";
    r41 := (r25 & r27 & r29 & r31 & r33 & r35 & r37 & r39);
    r43 := "1";
    r45 := "1";
    r47 := "1";
    r49 := "1";
    r51 := "1";
    r53 := "1";
    r55 := "1";
    r57 := "1";
    r59 := (r43 & r45 & r47 & r49 & r51 & r53 & r55 & r57);
    r61 := "1";
    r63 := "1";
    r65 := "1";
    r67 := "1";
    r69 := "1";
    r71 := "1";
    r73 := "1";
    r75 := "1";
    r77 := (r61 & r63 & r65 & r67 & r69 & r71 & r73 & r75);
    r79 := "1";
    r81 := "1";
    r83 := "1";
    r85 := "1";
    r87 := "1";
    r89 := "1";
    r91 := "1";
    r93 := "1";
    r95 := (r79 & r81 & r83 & r85 & r87 & r89 & r91 & r93);
    r97 := "1";
    r99 := "1";
    r101 := "1";
    r103 := "1";
    r105 := "1";
    r107 := "1";
    r109 := "1";
    r111 := "1";
    r113 := (r97 & r99 & r101 & r103 & r105 & r107 & r109 & r111);
    r115 := "1";
    r117 := "1";
    r119 := "1";
    r121 := "1";
    r123 := "1";
    r125 := "1";
    r127 := "1";
    r129 := "1";
    r131 := (r115 & r117 & r119 & r121 & r123 & r125 & r127 & r129);
    r133 := "1";
    r135 := "1";
    r137 := "1";
    r139 := "1";
    r141 := "1";
    r143 := "1";
    r145 := "1";
    r147 := "1";
    r149 := (r133 & r135 & r137 & r139 & r141 & r143 & r145 & r147);
    r151 := "1";
    r153 := "1";
    r155 := "1";
    r157 := "1";
    r159 := "1";
    r161 := "1";
    r163 := "1";
    r165 := "1";
    r167 := (r151 & r153 & r155 & r157 & r159 & r161 & r163 & r165);
    r169 := "1";
    r171 := "1";
    r173 := "1";
    r175 := "1";
    r177 := "1";
    r179 := "1";
    r181 := "1";
    r183 := "1";
    r185 := (r169 & r171 & r173 & r175 & r177 & r179 & r181 & r183);
    r187 := "1";
    r189 := "1";
    r191 := "1";
    r193 := "1";
    r195 := "1";
    r197 := "1";
    r199 := "1";
    r201 := "1";
    r203 := (r187 & r189 & r191 & r193 & r195 & r197 & r199 & r201);
    r205 := "1";
    r207 := "1";
    r209 := "1";
    r211 := "1";
    r213 := "1";
    r215 := "1";
    r217 := "1";
    r219 := "1";
    r221 := (r205 & r207 & r209 & r211 & r213 & r215 & r217 & r219);
    r223 := "1";
    r225 := "1";
    r227 := "1";
    r229 := "1";
    r231 := "1";
    r233 := "1";
    r235 := "1";
    r237 := "1";
    r239 := (r223 & r225 & r227 & r229 & r231 & r233 & r235 & r237);
    r241 := "1";
    r243 := "1";
    r245 := "1";
    r247 := "1";
    r249 := "1";
    r251 := "1";
    r253 := "1";
    r255 := "1";
    r257 := (r241 & r243 & r245 & r247 & r249 & r251 & r253 & r255);
    r259 := "1";
    r261 := "1";
    r263 := "1";
    r265 := "1";
    r267 := "1";
    r269 := "1";
    r271 := "1";
    r273 := "1";
    r275 := (r259 & r261 & r263 & r265 & r267 & r269 & r271 & r273);
    r277 := "1";
    r279 := "1";
    r281 := "1";
    r283 := "1";
    r285 := "1";
    r287 := "1";
    r289 := "1";
    r291 := "1";
    r293 := (r277 & r279 & r281 & r283 & r285 & r287 & r289 & r291);
    r295 := "1";
    r297 := "1";
    r299 := "1";
    r301 := "1";
    r303 := "1";
    r305 := "1";
    r307 := "1";
    r309 := "1";
    r311 := (r295 & r297 & r299 & r301 & r303 & r305 & r307 & r309);
    r313 := "1";
    r315 := "1";
    r317 := "1";
    r319 := "1";
    r321 := "1";
    r323 := "1";
    r325 := "1";
    r327 := "1";
    r329 := (r313 & r315 & r317 & r319 & r321 & r323 & r325 & r327);
    r331 := "1";
    r333 := "1";
    r335 := "1";
    r337 := "1";
    r339 := "1";
    r341 := "1";
    r343 := "1";
    r345 := "1";
    r347 := (r331 & r333 & r335 & r337 & r339 & r341 & r343 & r345);
    r349 := "1";
    r351 := "1";
    r353 := "1";
    r355 := "1";
    r357 := "1";
    r359 := "1";
    r361 := "1";
    r363 := "1";
    r365 := (r349 & r351 & r353 & r355 & r357 & r359 & r361 & r363);
    r367 := "1";
    r369 := "1";
    r371 := "1";
    r373 := "1";
    r375 := "1";
    r377 := "1";
    r379 := "1";
    r381 := "1";
    r383 := (r367 & r369 & r371 & r373 & r375 & r377 & r379 & r381);
    r385 := "1";
    r387 := "1";
    r389 := "1";
    r391 := "1";
    r393 := "1";
    r395 := "1";
    r397 := "1";
    r399 := "1";
    r401 := (r385 & r387 & r389 & r391 & r393 & r395 & r397 & r399);
    r403 := "1";
    r405 := "1";
    r407 := "1";
    r409 := "1";
    r411 := "1";
    r413 := "1";
    r415 := "1";
    r417 := "1";
    r419 := (r403 & r405 & r407 & r409 & r411 & r413 & r415 & r417);
    r421 := "1";
    r423 := "1";
    r425 := "1";
    r427 := "1";
    r429 := "1";
    r431 := "1";
    r433 := "1";
    r435 := "1";
    r437 := (r421 & r423 & r425 & r427 & r429 & r431 & r433 & r435);
    r439 := "1";
    r441 := "1";
    r443 := "1";
    r445 := "1";
    r447 := "1";
    r449 := "1";
    r451 := "1";
    r453 := "1";
    r455 := (r439 & r441 & r443 & r445 & r447 & r449 & r451 & r453);
    r457 := "1";
    r459 := "1";
    r461 := "1";
    r463 := "1";
    r465 := "1";
    r467 := "1";
    r469 := "1";
    r471 := "1";
    r473 := (r457 & r459 & r461 & r463 & r465 & r467 & r469 & r471);
    r475 := "1";
    r477 := "1";
    r479 := "1";
    r481 := "1";
    r483 := "1";
    r485 := "1";
    r487 := "1";
    r489 := "1";
    r491 := (r475 & r477 & r479 & r481 & r483 & r485 & r487 & r489);
    r493 := "1";
    r495 := "1";
    r497 := "1";
    r499 := "1";
    r501 := "1";
    r503 := "1";
    r505 := "1";
    r507 := "1";
    r509 := (r493 & r495 & r497 & r499 & r501 & r503 & r505 & r507);
    r511 := "1";
    r513 := "1";
    r515 := "1";
    r517 := "1";
    r519 := "1";
    r521 := "1";
    r523 := "1";
    r525 := "1";
    r527 := (r511 & r513 & r515 & r517 & r519 & r521 & r523 & r525);
    r529 := "1";
    r531 := "1";
    r533 := "1";
    r535 := "1";
    r537 := "1";
    r539 := "1";
    r541 := "1";
    r543 := "1";
    r545 := (r529 & r531 & r533 & r535 & r537 & r539 & r541 & r543);
    r547 := "1";
    r549 := "1";
    r551 := "1";
    r553 := "1";
    r555 := "1";
    r557 := "1";
    r559 := "1";
    r561 := "1";
    r563 := (r547 & r549 & r551 & r553 & r555 & r557 & r559 & r561);
    r565 := "1";
    r567 := "1";
    r569 := "1";
    r571 := "1";
    r573 := "1";
    r575 := "1";
    r577 := "1";
    r579 := "1";
    r581 := (r565 & r567 & r569 & r571 & r573 & r575 & r577 & r579);
    r583 := "1";
    r585 := "1";
    r587 := "1";
    r589 := "1";
    r591 := "1";
    r593 := "1";
    r595 := "1";
    r597 := "1";
    r599 := (r583 & r585 & r587 & r589 & r591 & r593 & r595 & r597);
    r601 := "1";
    r603 := "1";
    r605 := "1";
    r607 := "1";
    r609 := "1";
    r611 := "1";
    r613 := "1";
    r615 := "1";
    r617 := (r601 & r603 & r605 & r607 & r609 & r611 & r613 & r615);
    r619 := "1";
    r621 := "1";
    r623 := "1";
    r625 := "1";
    r627 := "1";
    r629 := "1";
    r631 := "1";
    r633 := "1";
    r635 := (r619 & r621 & r623 & r625 & r627 & r629 & r631 & r633);
    r637 := "1";
    r639 := "1";
    r641 := "1";
    r643 := "1";
    r645 := "1";
    r647 := "1";
    r649 := "1";
    r651 := "1";
    r653 := (r637 & r639 & r641 & r643 & r645 & r647 & r649 & r651);
    r655 := "1";
    r657 := "1";
    r659 := "1";
    r661 := "1";
    r663 := "1";
    r665 := "1";
    r667 := "1";
    r669 := "1";
    r671 := (r655 & r657 & r659 & r661 & r663 & r665 & r667 & r669);
    r673 := "1";
    r675 := "1";
    r677 := "1";
    r679 := "1";
    r681 := "1";
    r683 := "1";
    r685 := "1";
    r687 := "1";
    r689 := (r673 & r675 & r677 & r679 & r681 & r683 & r685 & r687);
    r691 := "1";
    r693 := "1";
    r695 := "1";
    r697 := "1";
    r699 := "1";
    r701 := "1";
    r703 := "1";
    r705 := "1";
    r707 := (r691 & r693 & r695 & r697 & r699 & r701 & r703 & r705);
    r709 := "1";
    r711 := "1";
    r713 := "1";
    r715 := "1";
    r717 := "1";
    r719 := "1";
    r721 := "1";
    r723 := "1";
    r725 := (r709 & r711 & r713 & r715 & r717 & r719 & r721 & r723);
    r727 := "1";
    r729 := "1";
    r731 := "1";
    r733 := "1";
    r735 := "1";
    r737 := "1";
    r739 := "1";
    r741 := "1";
    r743 := (r727 & r729 & r731 & r733 & r735 & r737 & r739 & r741);
    r745 := "1";
    r747 := "1";
    r749 := "1";
    r751 := "1";
    r753 := "1";
    r755 := "1";
    r757 := "1";
    r759 := "1";
    r761 := (r745 & r747 & r749 & r751 & r753 & r755 & r757 & r759);
    r763 := "1";
    r765 := "1";
    r767 := "1";
    r769 := "1";
    r771 := "1";
    r773 := "1";
    r775 := "1";
    r777 := "1";
    r779 := (r763 & r765 & r767 & r769 & r771 & r773 & r775 & r777);
    r781 := "1";
    r783 := "1";
    r785 := "1";
    r787 := "1";
    r789 := "1";
    r791 := "1";
    r793 := "1";
    r795 := "1";
    r797 := (r781 & r783 & r785 & r787 & r789 & r791 & r793 & r795);
    r799 := "1";
    r801 := "1";
    r803 := "1";
    r805 := "1";
    r807 := "1";
    r809 := "1";
    r811 := "1";
    r813 := "1";
    r815 := (r799 & r801 & r803 & r805 & r807 & r809 & r811 & r813);
    r817 := "1";
    r819 := "1";
    r821 := "1";
    r823 := "1";
    r825 := "1";
    r827 := "1";
    r829 := "1";
    r831 := "1";
    r833 := (r817 & r819 & r821 & r823 & r825 & r827 & r829 & r831);
    r835 := "1";
    r837 := "1";
    r839 := "1";
    r841 := "1";
    r843 := "1";
    r845 := "1";
    r847 := "1";
    r849 := "1";
    r851 := (r835 & r837 & r839 & r841 & r843 & r845 & r847 & r849);
    r853 := "1";
    r855 := "1";
    r857 := "1";
    r859 := "1";
    r861 := "1";
    r863 := "1";
    r865 := "1";
    r867 := "1";
    r869 := (r853 & r855 & r857 & r859 & r861 & r863 & r865 & r867);
    r871 := "1";
    r873 := "1";
    r875 := "1";
    r877 := "1";
    r879 := "1";
    r881 := "1";
    r883 := "1";
    r885 := "1";
    r887 := (r871 & r873 & r875 & r877 & r879 & r881 & r883 & r885);
    r889 := "1";
    r891 := "1";
    r893 := "1";
    r895 := "1";
    r897 := "1";
    r899 := "1";
    r901 := "1";
    r903 := "1";
    r905 := (r889 & r891 & r893 & r895 & r897 & r899 & r901 & r903);
    r907 := "1";
    r909 := "1";
    r911 := "1";
    r913 := "1";
    r915 := "1";
    r917 := "1";
    r919 := "1";
    r921 := "1";
    r923 := (r907 & r909 & r911 & r913 & r915 & r917 & r919 & r921);
    r925 := "1";
    r927 := "1";
    r929 := "1";
    r931 := "1";
    r933 := "1";
    r935 := "1";
    r937 := "1";
    r939 := "1";
    r941 := (r925 & r927 & r929 & r931 & r933 & r935 & r937 & r939);
    r943 := "1";
    r945 := "1";
    r947 := "1";
    r949 := "1";
    r951 := "1";
    r953 := "1";
    r955 := "1";
    r957 := "1";
    r959 := (r943 & r945 & r947 & r949 & r951 & r953 & r955 & r957);
    r961 := "1";
    r963 := "1";
    r965 := "1";
    r967 := "1";
    r969 := "1";
    r971 := "1";
    r973 := "1";
    r975 := "1";
    r977 := (r961 & r963 & r965 & r967 & r969 & r971 & r973 & r975);
    r979 := "1";
    r981 := "1";
    r983 := "1";
    r985 := "1";
    r987 := "1";
    r989 := "1";
    r991 := "1";
    r993 := "1";
    r995 := (r979 & r981 & r983 & r985 & r987 & r989 & r991 & r993);
    r997 := "1";
    r999 := "1";
    r1001 := "1";
    r1003 := "1";
    r1005 := "1";
    r1007 := "1";
    r1009 := "1";
    r1011 := "1";
    r1013 := (r997 & r999 & r1001 & r1003 & r1005 & r1007 & r1009 & r1011);
    r1015 := "1";
    r1017 := "1";
    r1019 := "1";
    r1021 := "1";
    r1023 := "1";
    r1025 := "1";
    r1027 := "1";
    r1029 := "1";
    r1031 := (r1015 & r1017 & r1019 & r1021 & r1023 & r1025 & r1027 & r1029);
    r1033 := "1";
    r1035 := "1";
    r1037 := "1";
    r1039 := "1";
    r1041 := "1";
    r1043 := "1";
    r1045 := "1";
    r1047 := "1";
    r1049 := (r1033 & r1035 & r1037 & r1039 & r1041 & r1043 & r1045 & r1047);
    r1051 := "1";
    r1053 := "1";
    r1055 := "1";
    r1057 := "1";
    r1059 := "1";
    r1061 := "1";
    r1063 := "1";
    r1065 := "1";
    r1067 := (r1051 & r1053 & r1055 & r1057 & r1059 & r1061 & r1063 & r1065);
    r1069 := "1";
    r1071 := "1";
    r1073 := "1";
    r1075 := "1";
    r1077 := "1";
    r1079 := "1";
    r1081 := "1";
    r1083 := "1";
    r1085 := (r1069 & r1071 & r1073 & r1075 & r1077 & r1079 & r1081 & r1083);
    r1087 := "1";
    r1089 := "1";
    r1091 := "1";
    r1093 := "1";
    r1095 := "1";
    r1097 := "1";
    r1099 := "1";
    r1101 := "1";
    r1103 := (r1087 & r1089 & r1091 & r1093 & r1095 & r1097 & r1099 & r1101);
    r1105 := "1";
    r1107 := "1";
    r1109 := "1";
    r1111 := "1";
    r1113 := "1";
    r1115 := "1";
    r1117 := "1";
    r1119 := "1";
    r1121 := (r1105 & r1107 & r1109 & r1111 & r1113 & r1115 & r1117 & r1119);
    r1123 := "1";
    r1125 := "1";
    r1127 := "1";
    r1129 := "1";
    r1131 := "1";
    r1133 := "1";
    r1135 := "1";
    r1137 := "1";
    r1139 := (r1123 & r1125 & r1127 & r1129 & r1131 & r1133 & r1135 & r1137);
    r1141 := "1";
    r1143 := "1";
    r1145 := "1";
    r1147 := "1";
    r1149 := "1";
    r1151 := "1";
    r1153 := "1";
    r1155 := "1";
    r1157 := (r1141 & r1143 & r1145 & r1147 & r1149 & r1151 & r1153 & r1155);
    r1158 := (r23 & r41 & r59 & r77 & r95 & r113 & r131 & r149 & r167 & r185 & r203 & r221 & r239 & r257 & r275 & r293 & r311 & r329 & r347 & r365 & r383 & r401 & r419 & r437 & r455 & r473 & r491 & r509 & r527 & r545 & r563 & r581 & r599 & r617 & r635 & r653 & r671 & r689 & r707 & r725 & r743 & r761 & r779 & r797 & r815 & r833 & r851 & r869 & r887 & r905 & r923 & r941 & r959 & r977 & r995 & r1013 & r1031 & r1049 & r1067 & r1085 & r1103 & r1121 & r1139 & r1157);
    return r1158;
  end rewire_zerothoutput_3;

begin
  process (clk)
    variable goto_L2965 : boolean := false;
    variable goto_L2959 : boolean := false;
    variable goto_L1163 : boolean := false;
    variable goto_L1165 : boolean := false;
    variable goto_L0 : boolean := false;
    variable goto_L2966 : boolean := false;
    variable r2958 : std_logic_vector(0 to 895) := (others => '0');
    variable r2955 : std_logic_vector(0 to 511) := (others => '0');
    variable r2951 : std_logic_vector(0 to 511) := (others => '0');
    variable r1195 : std_logic_vector(0 to 511) := (others => '0');
    variable r1194 : std_logic_vector(0 to 63) := (others => '0');
    variable r1193 : std_logic_vector(0 to 63) := (others => '0');
    variable r1192 : std_logic_vector(0 to 127) := (others => '0');
    variable r1191 : std_logic_vector(0 to 127) := (others => '0');
    variable b1188 : boolean := false;
    variable b1186 : boolean := false;
    variable b1184 : boolean := false;
    variable b1182 : boolean := false;
    variable b1180 : boolean := false;
    variable r1178 : std_logic_vector(0 to 511) := (others => '0');
    variable r1176 : std_logic_vector(0 to 63) := (others => '0');
    variable r1174 : std_logic_vector(0 to 63) := (others => '0');
    variable r1172 : std_logic_vector(0 to 127) := (others => '0');
    variable r1170 : std_logic_vector(0 to 127) := (others => '0');
    variable r1164 : std_logic_vector(0 to 895) := (others => '0');
    variable r1162 : std_logic_vector(0 to 895) := (others => '0');
    variable r1159 : std_logic_vector(0 to 511) := (others => '0');
    variable r4 : std_logic_vector(0 to 511) := (others => '0');
    variable state : control_state := STATE0;
  begin
    if clk'event and clk='1' then
      goto_L2965 := false;
      goto_L2959 := false;
      goto_L1163 := false;
      goto_L1165 := false;
      goto_L0 := false;
      goto_L2966 := false;
      null; -- label L2965
      -- ENTER
      goto_L0 := (state = STATE0);
      if (NOT goto_L0) then
        goto_L1163 := (state = STATE1163);
        if (NOT goto_L1163) then
          goto_L2959 := (state = STATE2959);
          null; -- label L2959
          r2958 := input;
          -- got r@J0 in r2958
          r1164 := r2958;
          goto_L1165 := true;
        end if;
        goto_L1165 := goto_L1165;
        if (NOT goto_L1165) then
          null; -- label L1163
          r1162 := input;
          -- got r@J1 in r1162
          r1164 := r1162;
          goto_L1165 := true;
        end if;
        goto_L1165 := goto_L1165;
        null; -- label L1165
        -- step in
        -- got x@IP in r1164
        -- final pat
        r1170 := r1164(0 to 127);
        r1172 := r1164(128 to 255);
        r1174 := r1164(256 to 319);
        r1176 := r1164(320 to 383);
        r1178 := r1164(384 to 895);
        b1180 := true;
        b1182 := true;
        b1184 := true;
        b1186 := true;
        b1188 := true;
        -- got key1@IQ in r1170
        -- got key2@IR in r1172
        -- got b0@IS in r1174
        -- got b1@IT in r1176
        r2951 := rewire_buildSalsa256_1190(r1170,r1172,r1174,r1176);
        -- got y@IV in r2951
        -- got b64@IU in r1178
        r2955 := xor512(r2951,r1178);
        output <= r2955;
        state := STATE2959;
        goto_L2966 := true;
      end if;
      goto_L2966 := goto_L2966;
      if (NOT goto_L2966) then
        null; -- label L0
        -- START
        -- foo in
        r1159 := rewire_zerothoutput_3;
        output <= r1159;
        state := STATE1163;
        goto_L2966 := true;
      end if;
      goto_L2966 := goto_L2966;
      null; -- label L2966
      -- EXIT
    end if;
  end process;
end behavioral;
library ieee;
use ieee.std_logic_1164.all;
-- Uncomment the following line if VHDL primitives are in use.
-- use prims.all;
entity main is
  Port ( clk : in std_logic ;
         input : in std_logic_vector (0 to 895);
         output : out std_logic_vector (0 to 511));
end main;
architecture structural of main is
begin
  dev : entity work.rwcomp0(behavioral)
    port map (clk,input,output);
    

end structural;
