library ieee;
use ieee.std_logic_1164.all;
-- Comment out the following line if VHDL primitives are not in use.
use work.prims.all;
entity rewire is
  Port ( clk : in std_logic ;
         input : in std_logic_vector (0 to 67);
         output : out std_logic_vector (0 to 64));
end rewire;

architecture behavioral of rewire is
  type control_state is (STATE0,STATE11,STATE686,STATE822,STATE958,STATE1094,STATE1230,STATE1366,STATE1502,STATE1638,STATE1784,STATE7570,STATE7728,STATE7767,STATE7806,STATE7844);
  function rewire_Maindigest3_7816(r7817 : std_logic_vector) return std_logic_vector;
  function rewire_Maindigest2_7778(r7779 : std_logic_vector) return std_logic_vector;
  function rewire_Maindigest1_7739(r7740 : std_logic_vector) return std_logic_vector;
  function rewire_Maindigest0_7700(r7701 : std_logic_vector) return std_logic_vector;
  function rewire_MainincCtr_7299(r7300 : std_logic_vector) return std_logic_vector;
  function rewire_Mainseed_2873(r2874 : std_logic_vector) return std_logic_vector;
  function rewire_MetaprogrammingRWwc67178f2_7224 return std_logic_vector;
  function rewire_MetaprogrammingRWwbef9a3f7_7155 return std_logic_vector;
  function rewire_MetaprogrammingRWwa4506ceb_7086 return std_logic_vector;
  function rewire_MetaprogrammingRWw90befffa_7017 return std_logic_vector;
  function rewire_MetaprogrammingRWw8cc70208_6948 return std_logic_vector;
  function rewire_MetaprogrammingRWw84c87814_6879 return std_logic_vector;
  function rewire_MetaprogrammingRWw78a5636f_6810 return std_logic_vector;
  function rewire_MetaprogrammingRWw748f82ee_6741 return std_logic_vector;
  function rewire_MetaprogrammingRWw682e6ff3_6672 return std_logic_vector;
  function rewire_MetaprogrammingRWw5b9cca4f_6603 return std_logic_vector;
  function rewire_MetaprogrammingRWw4ed8aa4a_6534 return std_logic_vector;
  function rewire_MetaprogrammingRWw391c0cb3_6465 return std_logic_vector;
  function rewire_MetaprogrammingRWw34b0bcb5_6396 return std_logic_vector;
  function rewire_MetaprogrammingRWw2748774c_6327 return std_logic_vector;
  function rewire_MetaprogrammingRWw1e376c08_6258 return std_logic_vector;
  function rewire_MetaprogrammingRWw19a4c116_6189 return std_logic_vector;
  function rewire_MetaprogrammingRWw106aa070_6120 return std_logic_vector;
  function rewire_MetaprogrammingRWwf40e3585_6051 return std_logic_vector;
  function rewire_MetaprogrammingRWwd6990624_5982 return std_logic_vector;
  function rewire_MetaprogrammingRWwd192e819_5913 return std_logic_vector;
  function rewire_MetaprogrammingRWwc76c51a3_5844 return std_logic_vector;
  function rewire_MetaprogrammingRWwc24b8b70_5775 return std_logic_vector;
  function rewire_MetaprogrammingRWwa81a664b_5706 return std_logic_vector;
  function rewire_MetaprogrammingRWwa2bfe8a1_5637 return std_logic_vector;
  function rewire_MetaprogrammingRWw92722c85_5568 return std_logic_vector;
  function rewire_MetaprogrammingRWw81c2c92e_5499 return std_logic_vector;
  function rewire_MetaprogrammingRWw766a0abb_5430 return std_logic_vector;
  function rewire_MetaprogrammingRWw650a7354_5361 return std_logic_vector;
  function rewire_MetaprogrammingRWw53380d13_5292 return std_logic_vector;
  function rewire_MetaprogrammingRWw4d2c6dfc_5223 return std_logic_vector;
  function rewire_MetaprogrammingRWw2e1b2138_5154 return std_logic_vector;
  function rewire_MetaprogrammingRWw27b70a85_5085 return std_logic_vector;
  function rewire_MetaprogrammingRWw14292967_5016 return std_logic_vector;
  function rewire_MetaprogrammingRWw06ca6351_4947 return std_logic_vector;
  function rewire_MetaprogrammingRWwd5a79147_4878 return std_logic_vector;
  function rewire_MetaprogrammingRWwc6e00bf3_4809 return std_logic_vector;
  function rewire_MetaprogrammingRWwbf597fc7_4740 return std_logic_vector;
  function rewire_MetaprogrammingRWwb00327c8_4671 return std_logic_vector;
  function rewire_MetaprogrammingRWwa831c66d_4602 return std_logic_vector;
  function rewire_MetaprogrammingRWw983e5152_4533 return std_logic_vector;
  function rewire_MetaprogrammingRWw76f988da_4464 return std_logic_vector;
  function rewire_MetaprogrammingRWw5cb0a9dc_4395 return std_logic_vector;
  function rewire_MetaprogrammingRWw4a7484aa_4326 return std_logic_vector;
  function rewire_MetaprogrammingRWw2de92c6f_4257 return std_logic_vector;
  function rewire_MetaprogrammingRWw240ca1cc_4188 return std_logic_vector;
  function rewire_MetaprogrammingRWw0fc19dc6_4119 return std_logic_vector;
  function rewire_MetaprogrammingRWwefbe4786_4050 return std_logic_vector;
  function rewire_MetaprogrammingRWwe49b69c1_3981 return std_logic_vector;
  function rewire_MetaprogrammingRWwc19bf174_3912 return std_logic_vector;
  function rewire_MetaprogrammingRWw9bdc06a7_3843 return std_logic_vector;
  function rewire_MetaprogrammingRWw80deb1fe_3774 return std_logic_vector;
  function rewire_MetaprogrammingRWw72be5d74_3705 return std_logic_vector;
  function rewire_MetaprogrammingRWw550c7dc3_3636 return std_logic_vector;
  function rewire_MetaprogrammingRWw243185be_3567 return std_logic_vector;
  function rewire_MetaprogrammingRWw12835b01_3498 return std_logic_vector;
  function rewire_MetaprogrammingRWwd807aa98_3429 return std_logic_vector;
  function rewire_MetaprogrammingRWwab1c5ed5_3360 return std_logic_vector;
  function rewire_MetaprogrammingRWw923f82a4_3291 return std_logic_vector;
  function rewire_MetaprogrammingRWw59f111f1_3222 return std_logic_vector;
  function rewire_MetaprogrammingRWw3956c25b_3153 return std_logic_vector;
  function rewire_MetaprogrammingRWwe9b5dba5_3084 return std_logic_vector;
  function rewire_MetaprogrammingRWwb5c0fbcf_3015 return std_logic_vector;
  function rewire_MetaprogrammingRWw71374491_2946 return std_logic_vector;
  function rewire_MetaprogrammingRWw428a2f98_2877 return std_logic_vector;
  function rewire_Mainstep256_2373(r2374 : std_logic_vector ; r2375 : std_logic_vector ; r2376 : std_logic_vector) return std_logic_vector;
  function rewire_Mainmaj_2854(r2855 : std_logic_vector ; r2856 : std_logic_vector ; r2857 : std_logic_vector) return std_logic_vector;
  function rewire_Mainbigsigma0_2636(r2637 : std_logic_vector) return std_logic_vector;
  function rewire_RWPreluderotateR22_2781(r2782 : std_logic_vector) return std_logic_vector;
  function rewire_RWPreluderotateR13_2709(r2710 : std_logic_vector) return std_logic_vector;
  function rewire_RWPreluderotateR2_2638(r2639 : std_logic_vector) return std_logic_vector;
  function rewire_Mainch_2623(r2624 : std_logic_vector ; r2625 : std_logic_vector ; r2626 : std_logic_vector) return std_logic_vector;
  function rewire_Mainbigsigma1_2405(r2406 : std_logic_vector) return std_logic_vector;
  function rewire_RWPreluderotateR25_2550(r2551 : std_logic_vector) return std_logic_vector;
  function rewire_RWPreluderotateR11_2478(r2479 : std_logic_vector) return std_logic_vector;
  function rewire_RWPreluderotateR6_2407(r2408 : std_logic_vector) return std_logic_vector;
  function rewire_MainupdateSched_1861(r1862 : std_logic_vector) return std_logic_vector;
  function rewire_Mainsigma0_2138(r2139 : std_logic_vector) return std_logic_vector;
  function rewire_RWPreludeshiftR3_2283(r2284 : std_logic_vector) return std_logic_vector;
  function rewire_RWPreluderotateR18_2211(r2212 : std_logic_vector) return std_logic_vector;
  function rewire_RWPreluderotateR7_2140(r2141 : std_logic_vector) return std_logic_vector;
  function rewire_Mainsigma1_1899(r1900 : std_logic_vector) return std_logic_vector;
  function rewire_RWPreludeshiftR10_2044(r2045 : std_logic_vector) return std_logic_vector;
  function rewire_RWPreluderotateR19_1972(r1973 : std_logic_vector) return std_logic_vector;
  function rewire_RWPreluderotateR17_1901(r1902 : std_logic_vector) return std_logic_vector;
  function rewire_MaininitialSHA256State_28 return std_logic_vector;
  function rewire_MetaprogrammingRWw5be0cd19_499 return std_logic_vector;
  function rewire_MetaprogrammingRWw1f83d9ab_432 return std_logic_vector;
  function rewire_MetaprogrammingRWw9b05688c_365 return std_logic_vector;
  function rewire_MetaprogrammingRWw510e527f_298 return std_logic_vector;
  function rewire_MetaprogrammingRWwa54ff53a_231 return std_logic_vector;
  function rewire_MetaprogrammingRWw3c6ef372_164 return std_logic_vector;
  function rewire_MetaprogrammingRWwbb67ae85_97 return std_logic_vector;
  function rewire_MetaprogrammingRWw6a09e667_30 return std_logic_vector;
  function rewire_Maindigest3_7816(r7817 : std_logic_vector) return std_logic_vector
  is
    variable r7838 : std_logic_vector(0 to 64) := (others => '0');
    variable r7837 : std_logic_vector(0 to 0) := (others => '0');
    variable b7836 : boolean := false;
    variable b7835 : boolean := false;
    variable b7834 : boolean := false;
    variable b7833 : boolean := false;
    variable b7832 : boolean := false;
    variable b7831 : boolean := false;
    variable b7830 : boolean := false;
    variable b7829 : boolean := false;
    variable b7828 : boolean := false;
    variable r7827 : std_logic_vector(0 to 31) := (others => '0');
    variable r7826 : std_logic_vector(0 to 31) := (others => '0');
    variable r7825 : std_logic_vector(0 to 31) := (others => '0');
    variable r7824 : std_logic_vector(0 to 31) := (others => '0');
    variable r7823 : std_logic_vector(0 to 31) := (others => '0');
    variable r7822 : std_logic_vector(0 to 31) := (others => '0');
    variable r7821 : std_logic_vector(0 to 31) := (others => '0');
    variable r7820 : std_logic_vector(0 to 31) := (others => '0');
    variable b7819 : boolean := false;
    variable r7818 : std_logic_vector(0 to 64) := (others => '0');
  begin
    null;
    b7819 := true;
    r7820 := r7817(0 to 31);
    r7821 := r7817(32 to 63);
    r7822 := r7817(64 to 95);
    r7823 := r7817(96 to 127);
    r7824 := r7817(128 to 159);
    r7825 := r7817(160 to 191);
    r7826 := r7817(192 to 223);
    r7827 := r7817(224 to 255);
    b7828 := true;
    b7829 := true;
    b7830 := true;
    b7831 := true;
    b7832 := true;
    b7833 := true;
    b7834 := true;
    b7835 := true;
    b7836 := (b7819 AND (b7828 AND (b7829 AND (b7830 AND (b7831 AND (b7832 AND (b7833 AND (b7834 AND b7835))))))));
    r7837 := "0";
    null;
    null;
    null;
    r7838 := (r7837 & r7826 & r7827);
    r7818 := r7838;
    return r7818;
  end rewire_Maindigest3_7816;
  function rewire_Maindigest2_7778(r7779 : std_logic_vector) return std_logic_vector
  is
    variable r7800 : std_logic_vector(0 to 64) := (others => '0');
    variable r7799 : std_logic_vector(0 to 0) := (others => '0');
    variable b7798 : boolean := false;
    variable b7797 : boolean := false;
    variable b7796 : boolean := false;
    variable b7795 : boolean := false;
    variable b7794 : boolean := false;
    variable b7793 : boolean := false;
    variable b7792 : boolean := false;
    variable b7791 : boolean := false;
    variable b7790 : boolean := false;
    variable r7789 : std_logic_vector(0 to 31) := (others => '0');
    variable r7788 : std_logic_vector(0 to 31) := (others => '0');
    variable r7787 : std_logic_vector(0 to 31) := (others => '0');
    variable r7786 : std_logic_vector(0 to 31) := (others => '0');
    variable r7785 : std_logic_vector(0 to 31) := (others => '0');
    variable r7784 : std_logic_vector(0 to 31) := (others => '0');
    variable r7783 : std_logic_vector(0 to 31) := (others => '0');
    variable r7782 : std_logic_vector(0 to 31) := (others => '0');
    variable b7781 : boolean := false;
    variable r7780 : std_logic_vector(0 to 64) := (others => '0');
  begin
    null;
    b7781 := true;
    r7782 := r7779(0 to 31);
    r7783 := r7779(32 to 63);
    r7784 := r7779(64 to 95);
    r7785 := r7779(96 to 127);
    r7786 := r7779(128 to 159);
    r7787 := r7779(160 to 191);
    r7788 := r7779(192 to 223);
    r7789 := r7779(224 to 255);
    b7790 := true;
    b7791 := true;
    b7792 := true;
    b7793 := true;
    b7794 := true;
    b7795 := true;
    b7796 := true;
    b7797 := true;
    b7798 := (b7781 AND (b7790 AND (b7791 AND (b7792 AND (b7793 AND (b7794 AND (b7795 AND (b7796 AND b7797))))))));
    r7799 := "0";
    null;
    null;
    null;
    r7800 := (r7799 & r7786 & r7787);
    r7780 := r7800;
    return r7780;
  end rewire_Maindigest2_7778;
  function rewire_Maindigest1_7739(r7740 : std_logic_vector) return std_logic_vector
  is
    variable r7761 : std_logic_vector(0 to 64) := (others => '0');
    variable r7760 : std_logic_vector(0 to 0) := (others => '0');
    variable b7759 : boolean := false;
    variable b7758 : boolean := false;
    variable b7757 : boolean := false;
    variable b7756 : boolean := false;
    variable b7755 : boolean := false;
    variable b7754 : boolean := false;
    variable b7753 : boolean := false;
    variable b7752 : boolean := false;
    variable b7751 : boolean := false;
    variable r7750 : std_logic_vector(0 to 31) := (others => '0');
    variable r7749 : std_logic_vector(0 to 31) := (others => '0');
    variable r7748 : std_logic_vector(0 to 31) := (others => '0');
    variable r7747 : std_logic_vector(0 to 31) := (others => '0');
    variable r7746 : std_logic_vector(0 to 31) := (others => '0');
    variable r7745 : std_logic_vector(0 to 31) := (others => '0');
    variable r7744 : std_logic_vector(0 to 31) := (others => '0');
    variable r7743 : std_logic_vector(0 to 31) := (others => '0');
    variable b7742 : boolean := false;
    variable r7741 : std_logic_vector(0 to 64) := (others => '0');
  begin
    null;
    b7742 := true;
    r7743 := r7740(0 to 31);
    r7744 := r7740(32 to 63);
    r7745 := r7740(64 to 95);
    r7746 := r7740(96 to 127);
    r7747 := r7740(128 to 159);
    r7748 := r7740(160 to 191);
    r7749 := r7740(192 to 223);
    r7750 := r7740(224 to 255);
    b7751 := true;
    b7752 := true;
    b7753 := true;
    b7754 := true;
    b7755 := true;
    b7756 := true;
    b7757 := true;
    b7758 := true;
    b7759 := (b7742 AND (b7751 AND (b7752 AND (b7753 AND (b7754 AND (b7755 AND (b7756 AND (b7757 AND b7758))))))));
    r7760 := "0";
    null;
    null;
    null;
    r7761 := (r7760 & r7745 & r7746);
    r7741 := r7761;
    return r7741;
  end rewire_Maindigest1_7739;
  function rewire_Maindigest0_7700(r7701 : std_logic_vector) return std_logic_vector
  is
    variable r7722 : std_logic_vector(0 to 64) := (others => '0');
    variable r7721 : std_logic_vector(0 to 0) := (others => '0');
    variable b7720 : boolean := false;
    variable b7719 : boolean := false;
    variable b7718 : boolean := false;
    variable b7717 : boolean := false;
    variable b7716 : boolean := false;
    variable b7715 : boolean := false;
    variable b7714 : boolean := false;
    variable b7713 : boolean := false;
    variable b7712 : boolean := false;
    variable r7711 : std_logic_vector(0 to 31) := (others => '0');
    variable r7710 : std_logic_vector(0 to 31) := (others => '0');
    variable r7709 : std_logic_vector(0 to 31) := (others => '0');
    variable r7708 : std_logic_vector(0 to 31) := (others => '0');
    variable r7707 : std_logic_vector(0 to 31) := (others => '0');
    variable r7706 : std_logic_vector(0 to 31) := (others => '0');
    variable r7705 : std_logic_vector(0 to 31) := (others => '0');
    variable r7704 : std_logic_vector(0 to 31) := (others => '0');
    variable b7703 : boolean := false;
    variable r7702 : std_logic_vector(0 to 64) := (others => '0');
  begin
    null;
    b7703 := true;
    r7704 := r7701(0 to 31);
    r7705 := r7701(32 to 63);
    r7706 := r7701(64 to 95);
    r7707 := r7701(96 to 127);
    r7708 := r7701(128 to 159);
    r7709 := r7701(160 to 191);
    r7710 := r7701(192 to 223);
    r7711 := r7701(224 to 255);
    b7712 := true;
    b7713 := true;
    b7714 := true;
    b7715 := true;
    b7716 := true;
    b7717 := true;
    b7718 := true;
    b7719 := true;
    b7720 := (b7703 AND (b7712 AND (b7713 AND (b7714 AND (b7715 AND (b7716 AND (b7717 AND (b7718 AND b7719))))))));
    r7721 := "0";
    null;
    null;
    null;
    r7722 := (r7721 & r7704 & r7705);
    r7702 := r7722;
    return r7702;
  end rewire_Maindigest0_7700;
  function rewire_MainincCtr_7299(r7300 : std_logic_vector) return std_logic_vector
  is
    variable r7556 : std_logic_vector(0 to 5) := (others => '0');
    variable r7555 : std_logic_vector(0 to 5) := (others => '0');
    variable b7554 : boolean := false;
    variable r7553 : std_logic_vector(0 to 5) := (others => '0');
    variable r7552 : std_logic_vector(0 to 5) := (others => '0');
    variable r7551 : std_logic_vector(0 to 5) := (others => '0');
    variable b7550 : boolean := false;
    variable r7549 : std_logic_vector(0 to 5) := (others => '0');
    variable r7548 : std_logic_vector(0 to 5) := (others => '0');
    variable r7547 : std_logic_vector(0 to 5) := (others => '0');
    variable b7546 : boolean := false;
    variable r7545 : std_logic_vector(0 to 5) := (others => '0');
    variable r7544 : std_logic_vector(0 to 5) := (others => '0');
    variable r7543 : std_logic_vector(0 to 5) := (others => '0');
    variable b7542 : boolean := false;
    variable r7541 : std_logic_vector(0 to 5) := (others => '0');
    variable r7540 : std_logic_vector(0 to 5) := (others => '0');
    variable r7539 : std_logic_vector(0 to 5) := (others => '0');
    variable b7538 : boolean := false;
    variable r7537 : std_logic_vector(0 to 5) := (others => '0');
    variable r7536 : std_logic_vector(0 to 5) := (others => '0');
    variable r7535 : std_logic_vector(0 to 5) := (others => '0');
    variable b7534 : boolean := false;
    variable r7533 : std_logic_vector(0 to 5) := (others => '0');
    variable r7532 : std_logic_vector(0 to 5) := (others => '0');
    variable r7531 : std_logic_vector(0 to 5) := (others => '0');
    variable b7530 : boolean := false;
    variable r7529 : std_logic_vector(0 to 5) := (others => '0');
    variable r7528 : std_logic_vector(0 to 5) := (others => '0');
    variable r7527 : std_logic_vector(0 to 5) := (others => '0');
    variable b7526 : boolean := false;
    variable r7525 : std_logic_vector(0 to 5) := (others => '0');
    variable r7524 : std_logic_vector(0 to 5) := (others => '0');
    variable r7523 : std_logic_vector(0 to 5) := (others => '0');
    variable b7522 : boolean := false;
    variable r7521 : std_logic_vector(0 to 5) := (others => '0');
    variable r7520 : std_logic_vector(0 to 5) := (others => '0');
    variable r7519 : std_logic_vector(0 to 5) := (others => '0');
    variable b7518 : boolean := false;
    variable r7517 : std_logic_vector(0 to 5) := (others => '0');
    variable r7516 : std_logic_vector(0 to 5) := (others => '0');
    variable r7515 : std_logic_vector(0 to 5) := (others => '0');
    variable b7514 : boolean := false;
    variable r7513 : std_logic_vector(0 to 5) := (others => '0');
    variable r7512 : std_logic_vector(0 to 5) := (others => '0');
    variable r7511 : std_logic_vector(0 to 5) := (others => '0');
    variable b7510 : boolean := false;
    variable r7509 : std_logic_vector(0 to 5) := (others => '0');
    variable r7508 : std_logic_vector(0 to 5) := (others => '0');
    variable r7507 : std_logic_vector(0 to 5) := (others => '0');
    variable b7506 : boolean := false;
    variable r7505 : std_logic_vector(0 to 5) := (others => '0');
    variable r7504 : std_logic_vector(0 to 5) := (others => '0');
    variable r7503 : std_logic_vector(0 to 5) := (others => '0');
    variable b7502 : boolean := false;
    variable r7501 : std_logic_vector(0 to 5) := (others => '0');
    variable r7500 : std_logic_vector(0 to 5) := (others => '0');
    variable r7499 : std_logic_vector(0 to 5) := (others => '0');
    variable b7498 : boolean := false;
    variable r7497 : std_logic_vector(0 to 5) := (others => '0');
    variable r7496 : std_logic_vector(0 to 5) := (others => '0');
    variable r7495 : std_logic_vector(0 to 5) := (others => '0');
    variable b7494 : boolean := false;
    variable r7493 : std_logic_vector(0 to 5) := (others => '0');
    variable r7492 : std_logic_vector(0 to 5) := (others => '0');
    variable r7491 : std_logic_vector(0 to 5) := (others => '0');
    variable b7490 : boolean := false;
    variable r7489 : std_logic_vector(0 to 5) := (others => '0');
    variable r7488 : std_logic_vector(0 to 5) := (others => '0');
    variable r7487 : std_logic_vector(0 to 5) := (others => '0');
    variable b7486 : boolean := false;
    variable r7485 : std_logic_vector(0 to 5) := (others => '0');
    variable r7484 : std_logic_vector(0 to 5) := (others => '0');
    variable r7483 : std_logic_vector(0 to 5) := (others => '0');
    variable b7482 : boolean := false;
    variable r7481 : std_logic_vector(0 to 5) := (others => '0');
    variable r7480 : std_logic_vector(0 to 5) := (others => '0');
    variable r7479 : std_logic_vector(0 to 5) := (others => '0');
    variable b7478 : boolean := false;
    variable r7477 : std_logic_vector(0 to 5) := (others => '0');
    variable r7476 : std_logic_vector(0 to 5) := (others => '0');
    variable r7475 : std_logic_vector(0 to 5) := (others => '0');
    variable b7474 : boolean := false;
    variable r7473 : std_logic_vector(0 to 5) := (others => '0');
    variable r7472 : std_logic_vector(0 to 5) := (others => '0');
    variable r7471 : std_logic_vector(0 to 5) := (others => '0');
    variable b7470 : boolean := false;
    variable r7469 : std_logic_vector(0 to 5) := (others => '0');
    variable r7468 : std_logic_vector(0 to 5) := (others => '0');
    variable r7467 : std_logic_vector(0 to 5) := (others => '0');
    variable b7466 : boolean := false;
    variable r7465 : std_logic_vector(0 to 5) := (others => '0');
    variable r7464 : std_logic_vector(0 to 5) := (others => '0');
    variable r7463 : std_logic_vector(0 to 5) := (others => '0');
    variable b7462 : boolean := false;
    variable r7461 : std_logic_vector(0 to 5) := (others => '0');
    variable r7460 : std_logic_vector(0 to 5) := (others => '0');
    variable r7459 : std_logic_vector(0 to 5) := (others => '0');
    variable b7458 : boolean := false;
    variable r7457 : std_logic_vector(0 to 5) := (others => '0');
    variable r7456 : std_logic_vector(0 to 5) := (others => '0');
    variable r7455 : std_logic_vector(0 to 5) := (others => '0');
    variable b7454 : boolean := false;
    variable r7453 : std_logic_vector(0 to 5) := (others => '0');
    variable r7452 : std_logic_vector(0 to 5) := (others => '0');
    variable r7451 : std_logic_vector(0 to 5) := (others => '0');
    variable b7450 : boolean := false;
    variable r7449 : std_logic_vector(0 to 5) := (others => '0');
    variable r7448 : std_logic_vector(0 to 5) := (others => '0');
    variable r7447 : std_logic_vector(0 to 5) := (others => '0');
    variable b7446 : boolean := false;
    variable r7445 : std_logic_vector(0 to 5) := (others => '0');
    variable r7444 : std_logic_vector(0 to 5) := (others => '0');
    variable r7443 : std_logic_vector(0 to 5) := (others => '0');
    variable b7442 : boolean := false;
    variable r7441 : std_logic_vector(0 to 5) := (others => '0');
    variable r7440 : std_logic_vector(0 to 5) := (others => '0');
    variable r7439 : std_logic_vector(0 to 5) := (others => '0');
    variable b7438 : boolean := false;
    variable r7437 : std_logic_vector(0 to 5) := (others => '0');
    variable r7436 : std_logic_vector(0 to 5) := (others => '0');
    variable r7435 : std_logic_vector(0 to 5) := (others => '0');
    variable b7434 : boolean := false;
    variable r7433 : std_logic_vector(0 to 5) := (others => '0');
    variable r7432 : std_logic_vector(0 to 5) := (others => '0');
    variable r7431 : std_logic_vector(0 to 5) := (others => '0');
    variable b7430 : boolean := false;
    variable r7429 : std_logic_vector(0 to 5) := (others => '0');
    variable r7428 : std_logic_vector(0 to 5) := (others => '0');
    variable r7427 : std_logic_vector(0 to 5) := (others => '0');
    variable b7426 : boolean := false;
    variable r7425 : std_logic_vector(0 to 5) := (others => '0');
    variable r7424 : std_logic_vector(0 to 5) := (others => '0');
    variable r7423 : std_logic_vector(0 to 5) := (others => '0');
    variable b7422 : boolean := false;
    variable r7421 : std_logic_vector(0 to 5) := (others => '0');
    variable r7420 : std_logic_vector(0 to 5) := (others => '0');
    variable r7419 : std_logic_vector(0 to 5) := (others => '0');
    variable b7418 : boolean := false;
    variable r7417 : std_logic_vector(0 to 5) := (others => '0');
    variable r7416 : std_logic_vector(0 to 5) := (others => '0');
    variable r7415 : std_logic_vector(0 to 5) := (others => '0');
    variable b7414 : boolean := false;
    variable r7413 : std_logic_vector(0 to 5) := (others => '0');
    variable r7412 : std_logic_vector(0 to 5) := (others => '0');
    variable r7411 : std_logic_vector(0 to 5) := (others => '0');
    variable b7410 : boolean := false;
    variable r7409 : std_logic_vector(0 to 5) := (others => '0');
    variable r7408 : std_logic_vector(0 to 5) := (others => '0');
    variable r7407 : std_logic_vector(0 to 5) := (others => '0');
    variable b7406 : boolean := false;
    variable r7405 : std_logic_vector(0 to 5) := (others => '0');
    variable r7404 : std_logic_vector(0 to 5) := (others => '0');
    variable r7403 : std_logic_vector(0 to 5) := (others => '0');
    variable b7402 : boolean := false;
    variable r7401 : std_logic_vector(0 to 5) := (others => '0');
    variable r7400 : std_logic_vector(0 to 5) := (others => '0');
    variable r7399 : std_logic_vector(0 to 5) := (others => '0');
    variable b7398 : boolean := false;
    variable r7397 : std_logic_vector(0 to 5) := (others => '0');
    variable r7396 : std_logic_vector(0 to 5) := (others => '0');
    variable r7395 : std_logic_vector(0 to 5) := (others => '0');
    variable b7394 : boolean := false;
    variable r7393 : std_logic_vector(0 to 5) := (others => '0');
    variable r7392 : std_logic_vector(0 to 5) := (others => '0');
    variable r7391 : std_logic_vector(0 to 5) := (others => '0');
    variable b7390 : boolean := false;
    variable r7389 : std_logic_vector(0 to 5) := (others => '0');
    variable r7388 : std_logic_vector(0 to 5) := (others => '0');
    variable r7387 : std_logic_vector(0 to 5) := (others => '0');
    variable b7386 : boolean := false;
    variable r7385 : std_logic_vector(0 to 5) := (others => '0');
    variable r7384 : std_logic_vector(0 to 5) := (others => '0');
    variable r7383 : std_logic_vector(0 to 5) := (others => '0');
    variable b7382 : boolean := false;
    variable r7381 : std_logic_vector(0 to 5) := (others => '0');
    variable r7380 : std_logic_vector(0 to 5) := (others => '0');
    variable r7379 : std_logic_vector(0 to 5) := (others => '0');
    variable b7378 : boolean := false;
    variable r7377 : std_logic_vector(0 to 5) := (others => '0');
    variable r7376 : std_logic_vector(0 to 5) := (others => '0');
    variable r7375 : std_logic_vector(0 to 5) := (others => '0');
    variable b7374 : boolean := false;
    variable r7373 : std_logic_vector(0 to 5) := (others => '0');
    variable r7372 : std_logic_vector(0 to 5) := (others => '0');
    variable r7371 : std_logic_vector(0 to 5) := (others => '0');
    variable b7370 : boolean := false;
    variable r7369 : std_logic_vector(0 to 5) := (others => '0');
    variable r7368 : std_logic_vector(0 to 5) := (others => '0');
    variable r7367 : std_logic_vector(0 to 5) := (others => '0');
    variable b7366 : boolean := false;
    variable r7365 : std_logic_vector(0 to 5) := (others => '0');
    variable r7364 : std_logic_vector(0 to 5) := (others => '0');
    variable r7363 : std_logic_vector(0 to 5) := (others => '0');
    variable b7362 : boolean := false;
    variable r7361 : std_logic_vector(0 to 5) := (others => '0');
    variable r7360 : std_logic_vector(0 to 5) := (others => '0');
    variable r7359 : std_logic_vector(0 to 5) := (others => '0');
    variable b7358 : boolean := false;
    variable r7357 : std_logic_vector(0 to 5) := (others => '0');
    variable r7356 : std_logic_vector(0 to 5) := (others => '0');
    variable r7355 : std_logic_vector(0 to 5) := (others => '0');
    variable b7354 : boolean := false;
    variable r7353 : std_logic_vector(0 to 5) := (others => '0');
    variable r7352 : std_logic_vector(0 to 5) := (others => '0');
    variable r7351 : std_logic_vector(0 to 5) := (others => '0');
    variable b7350 : boolean := false;
    variable r7349 : std_logic_vector(0 to 5) := (others => '0');
    variable r7348 : std_logic_vector(0 to 5) := (others => '0');
    variable r7347 : std_logic_vector(0 to 5) := (others => '0');
    variable b7346 : boolean := false;
    variable r7345 : std_logic_vector(0 to 5) := (others => '0');
    variable r7344 : std_logic_vector(0 to 5) := (others => '0');
    variable r7343 : std_logic_vector(0 to 5) := (others => '0');
    variable b7342 : boolean := false;
    variable r7341 : std_logic_vector(0 to 5) := (others => '0');
    variable r7340 : std_logic_vector(0 to 5) := (others => '0');
    variable r7339 : std_logic_vector(0 to 5) := (others => '0');
    variable b7338 : boolean := false;
    variable r7337 : std_logic_vector(0 to 5) := (others => '0');
    variable r7336 : std_logic_vector(0 to 5) := (others => '0');
    variable r7335 : std_logic_vector(0 to 5) := (others => '0');
    variable b7334 : boolean := false;
    variable r7333 : std_logic_vector(0 to 5) := (others => '0');
    variable r7332 : std_logic_vector(0 to 5) := (others => '0');
    variable r7331 : std_logic_vector(0 to 5) := (others => '0');
    variable b7330 : boolean := false;
    variable r7329 : std_logic_vector(0 to 5) := (others => '0');
    variable r7328 : std_logic_vector(0 to 5) := (others => '0');
    variable r7327 : std_logic_vector(0 to 5) := (others => '0');
    variable b7326 : boolean := false;
    variable r7325 : std_logic_vector(0 to 5) := (others => '0');
    variable r7324 : std_logic_vector(0 to 5) := (others => '0');
    variable r7323 : std_logic_vector(0 to 5) := (others => '0');
    variable b7322 : boolean := false;
    variable r7321 : std_logic_vector(0 to 5) := (others => '0');
    variable r7320 : std_logic_vector(0 to 5) := (others => '0');
    variable r7319 : std_logic_vector(0 to 5) := (others => '0');
    variable b7318 : boolean := false;
    variable r7317 : std_logic_vector(0 to 5) := (others => '0');
    variable r7316 : std_logic_vector(0 to 5) := (others => '0');
    variable r7315 : std_logic_vector(0 to 5) := (others => '0');
    variable b7314 : boolean := false;
    variable r7313 : std_logic_vector(0 to 5) := (others => '0');
    variable r7312 : std_logic_vector(0 to 5) := (others => '0');
    variable r7311 : std_logic_vector(0 to 5) := (others => '0');
    variable b7310 : boolean := false;
    variable r7309 : std_logic_vector(0 to 5) := (others => '0');
    variable r7308 : std_logic_vector(0 to 5) := (others => '0');
    variable r7307 : std_logic_vector(0 to 5) := (others => '0');
    variable b7306 : boolean := false;
    variable r7305 : std_logic_vector(0 to 5) := (others => '0');
    variable r7304 : std_logic_vector(0 to 5) := (others => '0');
    variable r7303 : std_logic_vector(0 to 5) := (others => '0');
    variable b7302 : boolean := false;
    variable r7301 : std_logic_vector(0 to 5) := (others => '0');
  begin
    null;
    b7302 := ("000000" = r7300(0 to 5));
    if b7302 then
      r7303 := "000001";
      null;
      r7304 := (r7303);
      r7301 := r7304;
     else 
      null;
      b7306 := ("000001" = r7300(0 to 5));
      if b7306 then
        r7307 := "000010";
        null;
        r7308 := (r7307);
        r7305 := r7308;
       else 
        null;
        b7310 := ("000010" = r7300(0 to 5));
        if b7310 then
          r7311 := "000011";
          null;
          r7312 := (r7311);
          r7309 := r7312;
         else 
          null;
          b7314 := ("000011" = r7300(0 to 5));
          if b7314 then
            r7315 := "000100";
            null;
            r7316 := (r7315);
            r7313 := r7316;
           else 
            null;
            b7318 := ("000100" = r7300(0 to 5));
            if b7318 then
              r7319 := "000101";
              null;
              r7320 := (r7319);
              r7317 := r7320;
             else 
              null;
              b7322 := ("000101" = r7300(0 to 5));
              if b7322 then
                r7323 := "000110";
                null;
                r7324 := (r7323);
                r7321 := r7324;
               else 
                null;
                b7326 := ("000110" = r7300(0 to 5));
                if b7326 then
                  r7327 := "000111";
                  null;
                  r7328 := (r7327);
                  r7325 := r7328;
                 else 
                  null;
                  b7330 := ("000111" = r7300(0 to 5));
                  if b7330 then
                    r7331 := "001000";
                    null;
                    r7332 := (r7331);
                    r7329 := r7332;
                   else 
                    null;
                    b7334 := ("001000" = r7300(0 to 5));
                    if b7334 then
                      r7335 := "001001";
                      null;
                      r7336 := (r7335);
                      r7333 := r7336;
                     else 
                      null;
                      b7338 := ("001001" = r7300(0 to 5));
                      if b7338 then
                        r7339 := "001010";
                        null;
                        r7340 := (r7339);
                        r7337 := r7340;
                       else 
                        null;
                        b7342 := ("001010" = r7300(0 to 5));
                        if b7342 then
                          r7343 := "001011";
                          null;
                          r7344 := (r7343);
                          r7341 := r7344;
                         else 
                          null;
                          b7346 := ("001011" = r7300(0 to 5));
                          if b7346 then
                            r7347 := "001100";
                            null;
                            r7348 := (r7347);
                            r7345 := r7348;
                           else 
                            null;
                            b7350 := ("001100" = r7300(0 to 5));
                            if b7350 then
                              r7351 := "001101";
                              null;
                              r7352 := (r7351);
                              r7349 := r7352;
                             else 
                              null;
                              b7354 := ("001101" = r7300(0 to 5));
                              if b7354 then
                                r7355 := "001110";
                                null;
                                r7356 := (r7355);
                                r7353 := r7356;
                               else 
                                null;
                                b7358 := ("001110" = r7300(0 to 5));
                                if b7358 then
                                  r7359 := "001111";
                                  null;
                                  r7360 := (r7359);
                                  r7357 := r7360;
                                 else 
                                  null;
                                  b7362 := ("001111" = r7300(0 to 5));
                                  if b7362 then
                                    r7363 := "010000";
                                    null;
                                    r7364 := (r7363);
                                    r7361 := r7364;
                                   else 
                                    null;
                                    b7366 := ("010000" = r7300(0 to 5));
                                    if b7366 then
                                      r7367 := "010001";
                                      null;
                                      r7368 := (r7367);
                                      r7365 := r7368;
                                     else 
                                      null;
                                      b7370 := ("010001" = r7300(0 to 5));
                                      if b7370 then
                                        r7371 := "010010";
                                        null;
                                        r7372 := (r7371);
                                        r7369 := r7372;
                                       else 
                                        null;
                                        b7374 := ("010010" = r7300(0 to 5));
                                        if b7374 then
                                          r7375 := "010011";
                                          null;
                                          r7376 := (r7375);
                                          r7373 := r7376;
                                         else 
                                          null;
                                          b7378 := ("010011" = r7300(0 to 5));
                                          if b7378 then
                                            r7379 := "010100";
                                            null;
                                            r7380 := (r7379);
                                            r7377 := r7380;
                                           else 
                                            null;
                                            b7382 := ("010100" = r7300(0 to 5));
                                            if b7382 then
                                              r7383 := "010101";
                                              null;
                                              r7384 := (r7383);
                                              r7381 := r7384;
                                             else 
                                              null;
                                              b7386 := ("010101" = r7300(0 to 5));
                                              if b7386 then
                                                r7387 := "010110";
                                                null;
                                                r7388 := (r7387);
                                                r7385 := r7388;
                                               else 
                                                null;
                                                b7390 := ("010110" = r7300(0 to 5));
                                                if b7390 then
                                                  r7391 := "010111";
                                                  null;
                                                  r7392 := (r7391);
                                                  r7389 := r7392;
                                                 else 
                                                  null;
                                                  b7394 := ("010111" = r7300(0 to 5));
                                                  if b7394 then
                                                    r7395 := "011000";
                                                    null;
                                                    r7396 := (r7395);
                                                    r7393 := r7396;
                                                   else 
                                                    null;
                                                    b7398 := ("011000" = r7300(0 to 5));
                                                    if b7398 then
                                                      r7399 := "011001";
                                                      null;
                                                      r7400 := (r7399);
                                                      r7397 := r7400;
                                                     else 
                                                      null;
                                                      b7402 := ("011001" = r7300(0 to 5));
                                                      if b7402 then
                                                        r7403 := "011010";
                                                        null;
                                                        r7404 := (r7403);
                                                        r7401 := r7404;
                                                       else 
                                                        null;
                                                        b7406 := ("011010" = r7300(0 to 5));
                                                        if b7406 then
                                                          r7407 := "011011";
                                                          null;
                                                          r7408 := (r7407);
                                                          r7405 := r7408;
                                                         else 
                                                          null;
                                                          b7410 := ("011011" = r7300(0 to 5));
                                                          if b7410 then
                                                            r7411 := "011100";
                                                            null;
                                                            r7412 := (r7411);
                                                            r7409 := r7412;
                                                           else 
                                                            null;
                                                            b7414 := ("011100" = r7300(0 to 5));
                                                            if b7414 then
                                                              r7415 := "011101";
                                                              null;
                                                              r7416 := (r7415);
                                                              r7413 := r7416;
                                                             else 
                                                              null;
                                                              b7418 := ("011101" = r7300(0 to 5));
                                                              if b7418 then
                                                                r7419 := "011110";
                                                                null;
                                                                r7420 := (r7419);
                                                                r7417 := r7420;
                                                               else 
                                                                null;
                                                                b7422 := ("011110" = r7300(0 to 5));
                                                                if b7422 then
                                                                  r7423 := "011111";
                                                                  null;
                                                                  r7424 := (r7423);
                                                                  r7421 := r7424;
                                                                 else 
                                                                  null;
                                                                  b7426 := ("011111" = r7300(0 to 5));
                                                                  if b7426 then
                                                                    r7427 := "100000";
                                                                    null;
                                                                    r7428 := (r7427);
                                                                    r7425 := r7428;
                                                                   else 
                                                                    null;
                                                                    b7430 := ("100000" = r7300(0 to 5));
                                                                    if b7430 then
                                                                      r7431 := "100001";
                                                                      null;
                                                                      r7432 := (r7431);
                                                                      r7429 := r7432;
                                                                     else 
                                                                      null;
                                                                      b7434 := ("100001" = r7300(0 to 5));
                                                                      if b7434 then
                                                                        r7435 := "100010";
                                                                        null;
                                                                        r7436 := (r7435);
                                                                        r7433 := r7436;
                                                                       else 
                                                                        null;
                                                                        b7438 := ("100010" = r7300(0 to 5));
                                                                        if b7438 then
                                                                          r7439 := "100011";
                                                                          null;
                                                                          r7440 := (r7439);
                                                                          r7437 := r7440;
                                                                         else 
                                                                          null;
                                                                          b7442 := ("100011" = r7300(0 to 5));
                                                                          if b7442 then
                                                                            r7443 := "100100";
                                                                            null;
                                                                            r7444 := (r7443);
                                                                            r7441 := r7444;
                                                                           else 
                                                                            null;
                                                                            b7446 := ("100100" = r7300(0 to 5));
                                                                            if b7446 then
                                                                              r7447 := "100101";
                                                                              null;
                                                                              r7448 := (r7447);
                                                                              r7445 := r7448;
                                                                             else 
                                                                              null;
                                                                              b7450 := ("100101" = r7300(0 to 5));
                                                                              if b7450 then
                                                                                r7451 := "100110";
                                                                                null;
                                                                                r7452 := (r7451);
                                                                                r7449 := r7452;
                                                                               else 
                                                                                null;
                                                                                b7454 := ("100110" = r7300(0 to 5));
                                                                                if b7454 then
                                                                                  r7455 := "100111";
                                                                                  null;
                                                                                  r7456 := (r7455);
                                                                                  r7453 := r7456;
                                                                                 else 
                                                                                  null;
                                                                                  b7458 := ("100111" = r7300(0 to 5));
                                                                                  if b7458 then
                                                                                    r7459 := "101000";
                                                                                    null;
                                                                                    r7460 := (r7459);
                                                                                    r7457 := r7460;
                                                                                   else 
                                                                                    null;
                                                                                    b7462 := ("101000" = r7300(0 to 5));
                                                                                    if b7462 then
                                                                                      r7463 := "101001";
                                                                                      null;
                                                                                      r7464 := (r7463);
                                                                                      r7461 := r7464;
                                                                                     else 
                                                                                      null;
                                                                                      b7466 := ("101001" = r7300(0 to 5));
                                                                                      if b7466 then
                                                                                        r7467 := "101010";
                                                                                        null;
                                                                                        r7468 := (r7467);
                                                                                        r7465 := r7468;
                                                                                       else 
                                                                                        null;
                                                                                        b7470 := ("101010" = r7300(0 to 5));
                                                                                        if b7470 then
                                                                                          r7471 := "101011";
                                                                                          null;
                                                                                          r7472 := (r7471);
                                                                                          r7469 := r7472;
                                                                                         else 
                                                                                          null;
                                                                                          b7474 := ("101011" = r7300(0 to 5));
                                                                                          if b7474 then
                                                                                            r7475 := "101100";
                                                                                            null;
                                                                                            r7476 := (r7475);
                                                                                            r7473 := r7476;
                                                                                           else 
                                                                                            null;
                                                                                            b7478 := ("101100" = r7300(0 to 5));
                                                                                            if b7478 then
                                                                                              r7479 := "101101";
                                                                                              null;
                                                                                              r7480 := (r7479);
                                                                                              r7477 := r7480;
                                                                                             else 
                                                                                              null;
                                                                                              b7482 := ("101101" = r7300(0 to 5));
                                                                                              if b7482 then
                                                                                                r7483 := "101110";
                                                                                                null;
                                                                                                r7484 := (r7483);
                                                                                                r7481 := r7484;
                                                                                               else 
                                                                                                null;
                                                                                                b7486 := ("101110" = r7300(0 to 5));
                                                                                                if b7486 then
                                                                                                  r7487 := "101111";
                                                                                                  null;
                                                                                                  r7488 := (r7487);
                                                                                                  r7485 := r7488;
                                                                                                 else 
                                                                                                  null;
                                                                                                  b7490 := ("101111" = r7300(0 to 5));
                                                                                                  if b7490 then
                                                                                                    r7491 := "110000";
                                                                                                    null;
                                                                                                    r7492 := (r7491);
                                                                                                    r7489 := r7492;
                                                                                                   else 
                                                                                                    null;
                                                                                                    b7494 := ("110000" = r7300(0 to 5));
                                                                                                    if b7494 then
                                                                                                      r7495 := "110001";
                                                                                                      null;
                                                                                                      r7496 := (r7495);
                                                                                                      r7493 := r7496;
                                                                                                     else 
                                                                                                      null;
                                                                                                      b7498 := ("110001" = r7300(0 to 5));
                                                                                                      if b7498 then
                                                                                                        r7499 := "110010";
                                                                                                        null;
                                                                                                        r7500 := (r7499);
                                                                                                        r7497 := r7500;
                                                                                                       else 
                                                                                                        null;
                                                                                                        b7502 := ("110010" = r7300(0 to 5));
                                                                                                        if b7502 then
                                                                                                          r7503 := "110011";
                                                                                                          null;
                                                                                                          r7504 := (r7503);
                                                                                                          r7501 := r7504;
                                                                                                         else 
                                                                                                          null;
                                                                                                          b7506 := ("110011" = r7300(0 to 5));
                                                                                                          if b7506 then
                                                                                                            r7507 := "110100";
                                                                                                            null;
                                                                                                            r7508 := (r7507);
                                                                                                            r7505 := r7508;
                                                                                                           else 
                                                                                                            null;
                                                                                                            b7510 := ("110100" = r7300(0 to 5));
                                                                                                            if b7510 then
                                                                                                              r7511 := "110101";
                                                                                                              null;
                                                                                                              r7512 := (r7511);
                                                                                                              r7509 := r7512;
                                                                                                             else 
                                                                                                              null;
                                                                                                              b7514 := ("110101" = r7300(0 to 5));
                                                                                                              if b7514 then
                                                                                                                r7515 := "110110";
                                                                                                                null;
                                                                                                                r7516 := (r7515);
                                                                                                                r7513 := r7516;
                                                                                                               else 
                                                                                                                null;
                                                                                                                b7518 := ("110110" = r7300(0 to 5));
                                                                                                                if b7518 then
                                                                                                                  r7519 := "110111";
                                                                                                                  null;
                                                                                                                  r7520 := (r7519);
                                                                                                                  r7517 := r7520;
                                                                                                                 else 
                                                                                                                  null;
                                                                                                                  b7522 := ("110111" = r7300(0 to 5));
                                                                                                                  if b7522 then
                                                                                                                    r7523 := "111000";
                                                                                                                    null;
                                                                                                                    r7524 := (r7523);
                                                                                                                    r7521 := r7524;
                                                                                                                   else 
                                                                                                                    null;
                                                                                                                    b7526 := ("111000" = r7300(0 to 5));
                                                                                                                    if b7526 then
                                                                                                                      r7527 := "111001";
                                                                                                                      null;
                                                                                                                      r7528 := (r7527);
                                                                                                                      r7525 := r7528;
                                                                                                                     else 
                                                                                                                      null;
                                                                                                                      b7530 := ("111001" = r7300(0 to 5));
                                                                                                                      if b7530 then
                                                                                                                        r7531 := "111010";
                                                                                                                        null;
                                                                                                                        r7532 := (r7531);
                                                                                                                        r7529 := r7532;
                                                                                                                       else 
                                                                                                                        null;
                                                                                                                        b7534 := ("111010" = r7300(0 to 5));
                                                                                                                        if b7534 then
                                                                                                                          r7535 := "111011";
                                                                                                                          null;
                                                                                                                          r7536 := (r7535);
                                                                                                                          r7533 := r7536;
                                                                                                                         else 
                                                                                                                          null;
                                                                                                                          b7538 := ("111011" = r7300(0 to 5));
                                                                                                                          if b7538 then
                                                                                                                            r7539 := "111100";
                                                                                                                            null;
                                                                                                                            r7540 := (r7539);
                                                                                                                            r7537 := r7540;
                                                                                                                           else 
                                                                                                                            null;
                                                                                                                            b7542 := ("111100" = r7300(0 to 5));
                                                                                                                            if b7542 then
                                                                                                                              r7543 := "111101";
                                                                                                                              null;
                                                                                                                              r7544 := (r7543);
                                                                                                                              r7541 := r7544;
                                                                                                                             else 
                                                                                                                              null;
                                                                                                                              b7546 := ("111101" = r7300(0 to 5));
                                                                                                                              if b7546 then
                                                                                                                                r7547 := "111110";
                                                                                                                                null;
                                                                                                                                r7548 := (r7547);
                                                                                                                                r7545 := r7548;
                                                                                                                               else 
                                                                                                                                null;
                                                                                                                                b7550 := ("111110" = r7300(0 to 5));
                                                                                                                                if b7550 then
                                                                                                                                  r7551 := "111111";
                                                                                                                                  null;
                                                                                                                                  r7552 := (r7551);
                                                                                                                                  r7549 := r7552;
                                                                                                                                 else 
                                                                                                                                  null;
                                                                                                                                  b7554 := ("111111" = r7300(0 to 5));
                                                                                                                                  r7555 := "000000";
                                                                                                                                  null;
                                                                                                                                  r7556 := (r7555);
                                                                                                                                  r7553 := r7556;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;
    return r7301;
  end rewire_MainincCtr_7299;
  function rewire_Mainseed_2873(r2874 : std_logic_vector) return std_logic_vector
  is
    variable r7290 : std_logic_vector(0 to 31) := (others => '0');
    variable b7223 : boolean := false;
    variable r7222 : std_logic_vector(0 to 31) := (others => '0');
    variable r7221 : std_logic_vector(0 to 31) := (others => '0');
    variable b7154 : boolean := false;
    variable r7153 : std_logic_vector(0 to 31) := (others => '0');
    variable r7152 : std_logic_vector(0 to 31) := (others => '0');
    variable b7085 : boolean := false;
    variable r7084 : std_logic_vector(0 to 31) := (others => '0');
    variable r7083 : std_logic_vector(0 to 31) := (others => '0');
    variable b7016 : boolean := false;
    variable r7015 : std_logic_vector(0 to 31) := (others => '0');
    variable r7014 : std_logic_vector(0 to 31) := (others => '0');
    variable b6947 : boolean := false;
    variable r6946 : std_logic_vector(0 to 31) := (others => '0');
    variable r6945 : std_logic_vector(0 to 31) := (others => '0');
    variable b6878 : boolean := false;
    variable r6877 : std_logic_vector(0 to 31) := (others => '0');
    variable r6876 : std_logic_vector(0 to 31) := (others => '0');
    variable b6809 : boolean := false;
    variable r6808 : std_logic_vector(0 to 31) := (others => '0');
    variable r6807 : std_logic_vector(0 to 31) := (others => '0');
    variable b6740 : boolean := false;
    variable r6739 : std_logic_vector(0 to 31) := (others => '0');
    variable r6738 : std_logic_vector(0 to 31) := (others => '0');
    variable b6671 : boolean := false;
    variable r6670 : std_logic_vector(0 to 31) := (others => '0');
    variable r6669 : std_logic_vector(0 to 31) := (others => '0');
    variable b6602 : boolean := false;
    variable r6601 : std_logic_vector(0 to 31) := (others => '0');
    variable r6600 : std_logic_vector(0 to 31) := (others => '0');
    variable b6533 : boolean := false;
    variable r6532 : std_logic_vector(0 to 31) := (others => '0');
    variable r6531 : std_logic_vector(0 to 31) := (others => '0');
    variable b6464 : boolean := false;
    variable r6463 : std_logic_vector(0 to 31) := (others => '0');
    variable r6462 : std_logic_vector(0 to 31) := (others => '0');
    variable b6395 : boolean := false;
    variable r6394 : std_logic_vector(0 to 31) := (others => '0');
    variable r6393 : std_logic_vector(0 to 31) := (others => '0');
    variable b6326 : boolean := false;
    variable r6325 : std_logic_vector(0 to 31) := (others => '0');
    variable r6324 : std_logic_vector(0 to 31) := (others => '0');
    variable b6257 : boolean := false;
    variable r6256 : std_logic_vector(0 to 31) := (others => '0');
    variable r6255 : std_logic_vector(0 to 31) := (others => '0');
    variable b6188 : boolean := false;
    variable r6187 : std_logic_vector(0 to 31) := (others => '0');
    variable r6186 : std_logic_vector(0 to 31) := (others => '0');
    variable b6119 : boolean := false;
    variable r6118 : std_logic_vector(0 to 31) := (others => '0');
    variable r6117 : std_logic_vector(0 to 31) := (others => '0');
    variable b6050 : boolean := false;
    variable r6049 : std_logic_vector(0 to 31) := (others => '0');
    variable r6048 : std_logic_vector(0 to 31) := (others => '0');
    variable b5981 : boolean := false;
    variable r5980 : std_logic_vector(0 to 31) := (others => '0');
    variable r5979 : std_logic_vector(0 to 31) := (others => '0');
    variable b5912 : boolean := false;
    variable r5911 : std_logic_vector(0 to 31) := (others => '0');
    variable r5910 : std_logic_vector(0 to 31) := (others => '0');
    variable b5843 : boolean := false;
    variable r5842 : std_logic_vector(0 to 31) := (others => '0');
    variable r5841 : std_logic_vector(0 to 31) := (others => '0');
    variable b5774 : boolean := false;
    variable r5773 : std_logic_vector(0 to 31) := (others => '0');
    variable r5772 : std_logic_vector(0 to 31) := (others => '0');
    variable b5705 : boolean := false;
    variable r5704 : std_logic_vector(0 to 31) := (others => '0');
    variable r5703 : std_logic_vector(0 to 31) := (others => '0');
    variable b5636 : boolean := false;
    variable r5635 : std_logic_vector(0 to 31) := (others => '0');
    variable r5634 : std_logic_vector(0 to 31) := (others => '0');
    variable b5567 : boolean := false;
    variable r5566 : std_logic_vector(0 to 31) := (others => '0');
    variable r5565 : std_logic_vector(0 to 31) := (others => '0');
    variable b5498 : boolean := false;
    variable r5497 : std_logic_vector(0 to 31) := (others => '0');
    variable r5496 : std_logic_vector(0 to 31) := (others => '0');
    variable b5429 : boolean := false;
    variable r5428 : std_logic_vector(0 to 31) := (others => '0');
    variable r5427 : std_logic_vector(0 to 31) := (others => '0');
    variable b5360 : boolean := false;
    variable r5359 : std_logic_vector(0 to 31) := (others => '0');
    variable r5358 : std_logic_vector(0 to 31) := (others => '0');
    variable b5291 : boolean := false;
    variable r5290 : std_logic_vector(0 to 31) := (others => '0');
    variable r5289 : std_logic_vector(0 to 31) := (others => '0');
    variable b5222 : boolean := false;
    variable r5221 : std_logic_vector(0 to 31) := (others => '0');
    variable r5220 : std_logic_vector(0 to 31) := (others => '0');
    variable b5153 : boolean := false;
    variable r5152 : std_logic_vector(0 to 31) := (others => '0');
    variable r5151 : std_logic_vector(0 to 31) := (others => '0');
    variable b5084 : boolean := false;
    variable r5083 : std_logic_vector(0 to 31) := (others => '0');
    variable r5082 : std_logic_vector(0 to 31) := (others => '0');
    variable b5015 : boolean := false;
    variable r5014 : std_logic_vector(0 to 31) := (others => '0');
    variable r5013 : std_logic_vector(0 to 31) := (others => '0');
    variable b4946 : boolean := false;
    variable r4945 : std_logic_vector(0 to 31) := (others => '0');
    variable r4944 : std_logic_vector(0 to 31) := (others => '0');
    variable b4877 : boolean := false;
    variable r4876 : std_logic_vector(0 to 31) := (others => '0');
    variable r4875 : std_logic_vector(0 to 31) := (others => '0');
    variable b4808 : boolean := false;
    variable r4807 : std_logic_vector(0 to 31) := (others => '0');
    variable r4806 : std_logic_vector(0 to 31) := (others => '0');
    variable b4739 : boolean := false;
    variable r4738 : std_logic_vector(0 to 31) := (others => '0');
    variable r4737 : std_logic_vector(0 to 31) := (others => '0');
    variable b4670 : boolean := false;
    variable r4669 : std_logic_vector(0 to 31) := (others => '0');
    variable r4668 : std_logic_vector(0 to 31) := (others => '0');
    variable b4601 : boolean := false;
    variable r4600 : std_logic_vector(0 to 31) := (others => '0');
    variable r4599 : std_logic_vector(0 to 31) := (others => '0');
    variable b4532 : boolean := false;
    variable r4531 : std_logic_vector(0 to 31) := (others => '0');
    variable r4530 : std_logic_vector(0 to 31) := (others => '0');
    variable b4463 : boolean := false;
    variable r4462 : std_logic_vector(0 to 31) := (others => '0');
    variable r4461 : std_logic_vector(0 to 31) := (others => '0');
    variable b4394 : boolean := false;
    variable r4393 : std_logic_vector(0 to 31) := (others => '0');
    variable r4392 : std_logic_vector(0 to 31) := (others => '0');
    variable b4325 : boolean := false;
    variable r4324 : std_logic_vector(0 to 31) := (others => '0');
    variable r4323 : std_logic_vector(0 to 31) := (others => '0');
    variable b4256 : boolean := false;
    variable r4255 : std_logic_vector(0 to 31) := (others => '0');
    variable r4254 : std_logic_vector(0 to 31) := (others => '0');
    variable b4187 : boolean := false;
    variable r4186 : std_logic_vector(0 to 31) := (others => '0');
    variable r4185 : std_logic_vector(0 to 31) := (others => '0');
    variable b4118 : boolean := false;
    variable r4117 : std_logic_vector(0 to 31) := (others => '0');
    variable r4116 : std_logic_vector(0 to 31) := (others => '0');
    variable b4049 : boolean := false;
    variable r4048 : std_logic_vector(0 to 31) := (others => '0');
    variable r4047 : std_logic_vector(0 to 31) := (others => '0');
    variable b3980 : boolean := false;
    variable r3979 : std_logic_vector(0 to 31) := (others => '0');
    variable r3978 : std_logic_vector(0 to 31) := (others => '0');
    variable b3911 : boolean := false;
    variable r3910 : std_logic_vector(0 to 31) := (others => '0');
    variable r3909 : std_logic_vector(0 to 31) := (others => '0');
    variable b3842 : boolean := false;
    variable r3841 : std_logic_vector(0 to 31) := (others => '0');
    variable r3840 : std_logic_vector(0 to 31) := (others => '0');
    variable b3773 : boolean := false;
    variable r3772 : std_logic_vector(0 to 31) := (others => '0');
    variable r3771 : std_logic_vector(0 to 31) := (others => '0');
    variable b3704 : boolean := false;
    variable r3703 : std_logic_vector(0 to 31) := (others => '0');
    variable r3702 : std_logic_vector(0 to 31) := (others => '0');
    variable b3635 : boolean := false;
    variable r3634 : std_logic_vector(0 to 31) := (others => '0');
    variable r3633 : std_logic_vector(0 to 31) := (others => '0');
    variable b3566 : boolean := false;
    variable r3565 : std_logic_vector(0 to 31) := (others => '0');
    variable r3564 : std_logic_vector(0 to 31) := (others => '0');
    variable b3497 : boolean := false;
    variable r3496 : std_logic_vector(0 to 31) := (others => '0');
    variable r3495 : std_logic_vector(0 to 31) := (others => '0');
    variable b3428 : boolean := false;
    variable r3427 : std_logic_vector(0 to 31) := (others => '0');
    variable r3426 : std_logic_vector(0 to 31) := (others => '0');
    variable b3359 : boolean := false;
    variable r3358 : std_logic_vector(0 to 31) := (others => '0');
    variable r3357 : std_logic_vector(0 to 31) := (others => '0');
    variable b3290 : boolean := false;
    variable r3289 : std_logic_vector(0 to 31) := (others => '0');
    variable r3288 : std_logic_vector(0 to 31) := (others => '0');
    variable b3221 : boolean := false;
    variable r3220 : std_logic_vector(0 to 31) := (others => '0');
    variable r3219 : std_logic_vector(0 to 31) := (others => '0');
    variable b3152 : boolean := false;
    variable r3151 : std_logic_vector(0 to 31) := (others => '0');
    variable r3150 : std_logic_vector(0 to 31) := (others => '0');
    variable b3083 : boolean := false;
    variable r3082 : std_logic_vector(0 to 31) := (others => '0');
    variable r3081 : std_logic_vector(0 to 31) := (others => '0');
    variable b3014 : boolean := false;
    variable r3013 : std_logic_vector(0 to 31) := (others => '0');
    variable r3012 : std_logic_vector(0 to 31) := (others => '0');
    variable b2945 : boolean := false;
    variable r2944 : std_logic_vector(0 to 31) := (others => '0');
    variable r2943 : std_logic_vector(0 to 31) := (others => '0');
    variable b2876 : boolean := false;
    variable r2875 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    b2876 := ("000000" = r2874(0 to 5));
    if b2876 then
      r2943 := rewire_MetaprogrammingRWw428a2f98_2877;
      r2875 := r2943;
     else 
      null;
      b2945 := ("000001" = r2874(0 to 5));
      if b2945 then
        r3012 := rewire_MetaprogrammingRWw71374491_2946;
        r2944 := r3012;
       else 
        null;
        b3014 := ("000010" = r2874(0 to 5));
        if b3014 then
          r3081 := rewire_MetaprogrammingRWwb5c0fbcf_3015;
          r3013 := r3081;
         else 
          null;
          b3083 := ("000011" = r2874(0 to 5));
          if b3083 then
            r3150 := rewire_MetaprogrammingRWwe9b5dba5_3084;
            r3082 := r3150;
           else 
            null;
            b3152 := ("000100" = r2874(0 to 5));
            if b3152 then
              r3219 := rewire_MetaprogrammingRWw3956c25b_3153;
              r3151 := r3219;
             else 
              null;
              b3221 := ("000101" = r2874(0 to 5));
              if b3221 then
                r3288 := rewire_MetaprogrammingRWw59f111f1_3222;
                r3220 := r3288;
               else 
                null;
                b3290 := ("000110" = r2874(0 to 5));
                if b3290 then
                  r3357 := rewire_MetaprogrammingRWw923f82a4_3291;
                  r3289 := r3357;
                 else 
                  null;
                  b3359 := ("000111" = r2874(0 to 5));
                  if b3359 then
                    r3426 := rewire_MetaprogrammingRWwab1c5ed5_3360;
                    r3358 := r3426;
                   else 
                    null;
                    b3428 := ("001000" = r2874(0 to 5));
                    if b3428 then
                      r3495 := rewire_MetaprogrammingRWwd807aa98_3429;
                      r3427 := r3495;
                     else 
                      null;
                      b3497 := ("001001" = r2874(0 to 5));
                      if b3497 then
                        r3564 := rewire_MetaprogrammingRWw12835b01_3498;
                        r3496 := r3564;
                       else 
                        null;
                        b3566 := ("001010" = r2874(0 to 5));
                        if b3566 then
                          r3633 := rewire_MetaprogrammingRWw243185be_3567;
                          r3565 := r3633;
                         else 
                          null;
                          b3635 := ("001011" = r2874(0 to 5));
                          if b3635 then
                            r3702 := rewire_MetaprogrammingRWw550c7dc3_3636;
                            r3634 := r3702;
                           else 
                            null;
                            b3704 := ("001100" = r2874(0 to 5));
                            if b3704 then
                              r3771 := rewire_MetaprogrammingRWw72be5d74_3705;
                              r3703 := r3771;
                             else 
                              null;
                              b3773 := ("001101" = r2874(0 to 5));
                              if b3773 then
                                r3840 := rewire_MetaprogrammingRWw80deb1fe_3774;
                                r3772 := r3840;
                               else 
                                null;
                                b3842 := ("001110" = r2874(0 to 5));
                                if b3842 then
                                  r3909 := rewire_MetaprogrammingRWw9bdc06a7_3843;
                                  r3841 := r3909;
                                 else 
                                  null;
                                  b3911 := ("001111" = r2874(0 to 5));
                                  if b3911 then
                                    r3978 := rewire_MetaprogrammingRWwc19bf174_3912;
                                    r3910 := r3978;
                                   else 
                                    null;
                                    b3980 := ("010000" = r2874(0 to 5));
                                    if b3980 then
                                      r4047 := rewire_MetaprogrammingRWwe49b69c1_3981;
                                      r3979 := r4047;
                                     else 
                                      null;
                                      b4049 := ("010001" = r2874(0 to 5));
                                      if b4049 then
                                        r4116 := rewire_MetaprogrammingRWwefbe4786_4050;
                                        r4048 := r4116;
                                       else 
                                        null;
                                        b4118 := ("010010" = r2874(0 to 5));
                                        if b4118 then
                                          r4185 := rewire_MetaprogrammingRWw0fc19dc6_4119;
                                          r4117 := r4185;
                                         else 
                                          null;
                                          b4187 := ("010011" = r2874(0 to 5));
                                          if b4187 then
                                            r4254 := rewire_MetaprogrammingRWw240ca1cc_4188;
                                            r4186 := r4254;
                                           else 
                                            null;
                                            b4256 := ("010100" = r2874(0 to 5));
                                            if b4256 then
                                              r4323 := rewire_MetaprogrammingRWw2de92c6f_4257;
                                              r4255 := r4323;
                                             else 
                                              null;
                                              b4325 := ("010101" = r2874(0 to 5));
                                              if b4325 then
                                                r4392 := rewire_MetaprogrammingRWw4a7484aa_4326;
                                                r4324 := r4392;
                                               else 
                                                null;
                                                b4394 := ("010110" = r2874(0 to 5));
                                                if b4394 then
                                                  r4461 := rewire_MetaprogrammingRWw5cb0a9dc_4395;
                                                  r4393 := r4461;
                                                 else 
                                                  null;
                                                  b4463 := ("010111" = r2874(0 to 5));
                                                  if b4463 then
                                                    r4530 := rewire_MetaprogrammingRWw76f988da_4464;
                                                    r4462 := r4530;
                                                   else 
                                                    null;
                                                    b4532 := ("011000" = r2874(0 to 5));
                                                    if b4532 then
                                                      r4599 := rewire_MetaprogrammingRWw983e5152_4533;
                                                      r4531 := r4599;
                                                     else 
                                                      null;
                                                      b4601 := ("011001" = r2874(0 to 5));
                                                      if b4601 then
                                                        r4668 := rewire_MetaprogrammingRWwa831c66d_4602;
                                                        r4600 := r4668;
                                                       else 
                                                        null;
                                                        b4670 := ("011010" = r2874(0 to 5));
                                                        if b4670 then
                                                          r4737 := rewire_MetaprogrammingRWwb00327c8_4671;
                                                          r4669 := r4737;
                                                         else 
                                                          null;
                                                          b4739 := ("011011" = r2874(0 to 5));
                                                          if b4739 then
                                                            r4806 := rewire_MetaprogrammingRWwbf597fc7_4740;
                                                            r4738 := r4806;
                                                           else 
                                                            null;
                                                            b4808 := ("011100" = r2874(0 to 5));
                                                            if b4808 then
                                                              r4875 := rewire_MetaprogrammingRWwc6e00bf3_4809;
                                                              r4807 := r4875;
                                                             else 
                                                              null;
                                                              b4877 := ("011101" = r2874(0 to 5));
                                                              if b4877 then
                                                                r4944 := rewire_MetaprogrammingRWwd5a79147_4878;
                                                                r4876 := r4944;
                                                               else 
                                                                null;
                                                                b4946 := ("011110" = r2874(0 to 5));
                                                                if b4946 then
                                                                  r5013 := rewire_MetaprogrammingRWw06ca6351_4947;
                                                                  r4945 := r5013;
                                                                 else 
                                                                  null;
                                                                  b5015 := ("011111" = r2874(0 to 5));
                                                                  if b5015 then
                                                                    r5082 := rewire_MetaprogrammingRWw14292967_5016;
                                                                    r5014 := r5082;
                                                                   else 
                                                                    null;
                                                                    b5084 := ("100000" = r2874(0 to 5));
                                                                    if b5084 then
                                                                      r5151 := rewire_MetaprogrammingRWw27b70a85_5085;
                                                                      r5083 := r5151;
                                                                     else 
                                                                      null;
                                                                      b5153 := ("100001" = r2874(0 to 5));
                                                                      if b5153 then
                                                                        r5220 := rewire_MetaprogrammingRWw2e1b2138_5154;
                                                                        r5152 := r5220;
                                                                       else 
                                                                        null;
                                                                        b5222 := ("100010" = r2874(0 to 5));
                                                                        if b5222 then
                                                                          r5289 := rewire_MetaprogrammingRWw4d2c6dfc_5223;
                                                                          r5221 := r5289;
                                                                         else 
                                                                          null;
                                                                          b5291 := ("100011" = r2874(0 to 5));
                                                                          if b5291 then
                                                                            r5358 := rewire_MetaprogrammingRWw53380d13_5292;
                                                                            r5290 := r5358;
                                                                           else 
                                                                            null;
                                                                            b5360 := ("100100" = r2874(0 to 5));
                                                                            if b5360 then
                                                                              r5427 := rewire_MetaprogrammingRWw650a7354_5361;
                                                                              r5359 := r5427;
                                                                             else 
                                                                              null;
                                                                              b5429 := ("100101" = r2874(0 to 5));
                                                                              if b5429 then
                                                                                r5496 := rewire_MetaprogrammingRWw766a0abb_5430;
                                                                                r5428 := r5496;
                                                                               else 
                                                                                null;
                                                                                b5498 := ("100110" = r2874(0 to 5));
                                                                                if b5498 then
                                                                                  r5565 := rewire_MetaprogrammingRWw81c2c92e_5499;
                                                                                  r5497 := r5565;
                                                                                 else 
                                                                                  null;
                                                                                  b5567 := ("100111" = r2874(0 to 5));
                                                                                  if b5567 then
                                                                                    r5634 := rewire_MetaprogrammingRWw92722c85_5568;
                                                                                    r5566 := r5634;
                                                                                   else 
                                                                                    null;
                                                                                    b5636 := ("101000" = r2874(0 to 5));
                                                                                    if b5636 then
                                                                                      r5703 := rewire_MetaprogrammingRWwa2bfe8a1_5637;
                                                                                      r5635 := r5703;
                                                                                     else 
                                                                                      null;
                                                                                      b5705 := ("101001" = r2874(0 to 5));
                                                                                      if b5705 then
                                                                                        r5772 := rewire_MetaprogrammingRWwa81a664b_5706;
                                                                                        r5704 := r5772;
                                                                                       else 
                                                                                        null;
                                                                                        b5774 := ("101010" = r2874(0 to 5));
                                                                                        if b5774 then
                                                                                          r5841 := rewire_MetaprogrammingRWwc24b8b70_5775;
                                                                                          r5773 := r5841;
                                                                                         else 
                                                                                          null;
                                                                                          b5843 := ("101011" = r2874(0 to 5));
                                                                                          if b5843 then
                                                                                            r5910 := rewire_MetaprogrammingRWwc76c51a3_5844;
                                                                                            r5842 := r5910;
                                                                                           else 
                                                                                            null;
                                                                                            b5912 := ("101100" = r2874(0 to 5));
                                                                                            if b5912 then
                                                                                              r5979 := rewire_MetaprogrammingRWwd192e819_5913;
                                                                                              r5911 := r5979;
                                                                                             else 
                                                                                              null;
                                                                                              b5981 := ("101101" = r2874(0 to 5));
                                                                                              if b5981 then
                                                                                                r6048 := rewire_MetaprogrammingRWwd6990624_5982;
                                                                                                r5980 := r6048;
                                                                                               else 
                                                                                                null;
                                                                                                b6050 := ("101110" = r2874(0 to 5));
                                                                                                if b6050 then
                                                                                                  r6117 := rewire_MetaprogrammingRWwf40e3585_6051;
                                                                                                  r6049 := r6117;
                                                                                                 else 
                                                                                                  null;
                                                                                                  b6119 := ("101111" = r2874(0 to 5));
                                                                                                  if b6119 then
                                                                                                    r6186 := rewire_MetaprogrammingRWw106aa070_6120;
                                                                                                    r6118 := r6186;
                                                                                                   else 
                                                                                                    null;
                                                                                                    b6188 := ("110000" = r2874(0 to 5));
                                                                                                    if b6188 then
                                                                                                      r6255 := rewire_MetaprogrammingRWw19a4c116_6189;
                                                                                                      r6187 := r6255;
                                                                                                     else 
                                                                                                      null;
                                                                                                      b6257 := ("110001" = r2874(0 to 5));
                                                                                                      if b6257 then
                                                                                                        r6324 := rewire_MetaprogrammingRWw1e376c08_6258;
                                                                                                        r6256 := r6324;
                                                                                                       else 
                                                                                                        null;
                                                                                                        b6326 := ("110010" = r2874(0 to 5));
                                                                                                        if b6326 then
                                                                                                          r6393 := rewire_MetaprogrammingRWw2748774c_6327;
                                                                                                          r6325 := r6393;
                                                                                                         else 
                                                                                                          null;
                                                                                                          b6395 := ("110011" = r2874(0 to 5));
                                                                                                          if b6395 then
                                                                                                            r6462 := rewire_MetaprogrammingRWw34b0bcb5_6396;
                                                                                                            r6394 := r6462;
                                                                                                           else 
                                                                                                            null;
                                                                                                            b6464 := ("110100" = r2874(0 to 5));
                                                                                                            if b6464 then
                                                                                                              r6531 := rewire_MetaprogrammingRWw391c0cb3_6465;
                                                                                                              r6463 := r6531;
                                                                                                             else 
                                                                                                              null;
                                                                                                              b6533 := ("110101" = r2874(0 to 5));
                                                                                                              if b6533 then
                                                                                                                r6600 := rewire_MetaprogrammingRWw4ed8aa4a_6534;
                                                                                                                r6532 := r6600;
                                                                                                               else 
                                                                                                                null;
                                                                                                                b6602 := ("110110" = r2874(0 to 5));
                                                                                                                if b6602 then
                                                                                                                  r6669 := rewire_MetaprogrammingRWw5b9cca4f_6603;
                                                                                                                  r6601 := r6669;
                                                                                                                 else 
                                                                                                                  null;
                                                                                                                  b6671 := ("110111" = r2874(0 to 5));
                                                                                                                  if b6671 then
                                                                                                                    r6738 := rewire_MetaprogrammingRWw682e6ff3_6672;
                                                                                                                    r6670 := r6738;
                                                                                                                   else 
                                                                                                                    null;
                                                                                                                    b6740 := ("111000" = r2874(0 to 5));
                                                                                                                    if b6740 then
                                                                                                                      r6807 := rewire_MetaprogrammingRWw748f82ee_6741;
                                                                                                                      r6739 := r6807;
                                                                                                                     else 
                                                                                                                      null;
                                                                                                                      b6809 := ("111001" = r2874(0 to 5));
                                                                                                                      if b6809 then
                                                                                                                        r6876 := rewire_MetaprogrammingRWw78a5636f_6810;
                                                                                                                        r6808 := r6876;
                                                                                                                       else 
                                                                                                                        null;
                                                                                                                        b6878 := ("111010" = r2874(0 to 5));
                                                                                                                        if b6878 then
                                                                                                                          r6945 := rewire_MetaprogrammingRWw84c87814_6879;
                                                                                                                          r6877 := r6945;
                                                                                                                         else 
                                                                                                                          null;
                                                                                                                          b6947 := ("111011" = r2874(0 to 5));
                                                                                                                          if b6947 then
                                                                                                                            r7014 := rewire_MetaprogrammingRWw8cc70208_6948;
                                                                                                                            r6946 := r7014;
                                                                                                                           else 
                                                                                                                            null;
                                                                                                                            b7016 := ("111100" = r2874(0 to 5));
                                                                                                                            if b7016 then
                                                                                                                              r7083 := rewire_MetaprogrammingRWw90befffa_7017;
                                                                                                                              r7015 := r7083;
                                                                                                                             else 
                                                                                                                              null;
                                                                                                                              b7085 := ("111101" = r2874(0 to 5));
                                                                                                                              if b7085 then
                                                                                                                                r7152 := rewire_MetaprogrammingRWwa4506ceb_7086;
                                                                                                                                r7084 := r7152;
                                                                                                                               else 
                                                                                                                                null;
                                                                                                                                b7154 := ("111110" = r2874(0 to 5));
                                                                                                                                if b7154 then
                                                                                                                                  r7221 := rewire_MetaprogrammingRWwbef9a3f7_7155;
                                                                                                                                  r7153 := r7221;
                                                                                                                                 else 
                                                                                                                                  null;
                                                                                                                                  b7223 := ("111111" = r2874(0 to 5));
                                                                                                                                  r7290 := rewire_MetaprogrammingRWwc67178f2_7224;
                                                                                                                                  r7222 := r7290;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;
    return r2875;
  end rewire_Mainseed_2873;
  function rewire_MetaprogrammingRWwc67178f2_7224 return std_logic_vector
  is
    variable r7289 : std_logic_vector(0 to 0) := (others => '0');
    variable r7288 : std_logic_vector(0 to 0) := (others => '0');
    variable r7287 : std_logic_vector(0 to 0) := (others => '0');
    variable r7286 : std_logic_vector(0 to 0) := (others => '0');
    variable r7285 : std_logic_vector(0 to 0) := (others => '0');
    variable r7284 : std_logic_vector(0 to 0) := (others => '0');
    variable r7283 : std_logic_vector(0 to 0) := (others => '0');
    variable r7282 : std_logic_vector(0 to 0) := (others => '0');
    variable r7281 : std_logic_vector(0 to 0) := (others => '0');
    variable r7280 : std_logic_vector(0 to 0) := (others => '0');
    variable r7279 : std_logic_vector(0 to 0) := (others => '0');
    variable r7278 : std_logic_vector(0 to 0) := (others => '0');
    variable r7277 : std_logic_vector(0 to 0) := (others => '0');
    variable r7276 : std_logic_vector(0 to 0) := (others => '0');
    variable r7275 : std_logic_vector(0 to 0) := (others => '0');
    variable r7274 : std_logic_vector(0 to 0) := (others => '0');
    variable r7273 : std_logic_vector(0 to 0) := (others => '0');
    variable r7272 : std_logic_vector(0 to 0) := (others => '0');
    variable r7271 : std_logic_vector(0 to 0) := (others => '0');
    variable r7270 : std_logic_vector(0 to 0) := (others => '0');
    variable r7269 : std_logic_vector(0 to 0) := (others => '0');
    variable r7268 : std_logic_vector(0 to 0) := (others => '0');
    variable r7267 : std_logic_vector(0 to 0) := (others => '0');
    variable r7266 : std_logic_vector(0 to 0) := (others => '0');
    variable r7265 : std_logic_vector(0 to 0) := (others => '0');
    variable r7264 : std_logic_vector(0 to 0) := (others => '0');
    variable r7263 : std_logic_vector(0 to 0) := (others => '0');
    variable r7262 : std_logic_vector(0 to 0) := (others => '0');
    variable r7261 : std_logic_vector(0 to 0) := (others => '0');
    variable r7260 : std_logic_vector(0 to 0) := (others => '0');
    variable r7259 : std_logic_vector(0 to 0) := (others => '0');
    variable r7258 : std_logic_vector(0 to 0) := (others => '0');
    variable r7257 : std_logic_vector(0 to 0) := (others => '0');
    variable r7256 : std_logic_vector(0 to 0) := (others => '0');
    variable r7255 : std_logic_vector(0 to 0) := (others => '0');
    variable r7254 : std_logic_vector(0 to 0) := (others => '0');
    variable r7253 : std_logic_vector(0 to 0) := (others => '0');
    variable r7252 : std_logic_vector(0 to 0) := (others => '0');
    variable r7251 : std_logic_vector(0 to 0) := (others => '0');
    variable r7250 : std_logic_vector(0 to 0) := (others => '0');
    variable r7249 : std_logic_vector(0 to 0) := (others => '0');
    variable r7248 : std_logic_vector(0 to 0) := (others => '0');
    variable r7247 : std_logic_vector(0 to 0) := (others => '0');
    variable r7246 : std_logic_vector(0 to 0) := (others => '0');
    variable r7245 : std_logic_vector(0 to 0) := (others => '0');
    variable r7244 : std_logic_vector(0 to 0) := (others => '0');
    variable r7243 : std_logic_vector(0 to 0) := (others => '0');
    variable r7242 : std_logic_vector(0 to 0) := (others => '0');
    variable r7241 : std_logic_vector(0 to 0) := (others => '0');
    variable r7240 : std_logic_vector(0 to 0) := (others => '0');
    variable r7239 : std_logic_vector(0 to 0) := (others => '0');
    variable r7238 : std_logic_vector(0 to 0) := (others => '0');
    variable r7237 : std_logic_vector(0 to 0) := (others => '0');
    variable r7236 : std_logic_vector(0 to 0) := (others => '0');
    variable r7235 : std_logic_vector(0 to 0) := (others => '0');
    variable r7234 : std_logic_vector(0 to 0) := (others => '0');
    variable r7233 : std_logic_vector(0 to 0) := (others => '0');
    variable r7232 : std_logic_vector(0 to 0) := (others => '0');
    variable r7231 : std_logic_vector(0 to 0) := (others => '0');
    variable r7230 : std_logic_vector(0 to 0) := (others => '0');
    variable r7229 : std_logic_vector(0 to 0) := (others => '0');
    variable r7228 : std_logic_vector(0 to 0) := (others => '0');
    variable r7227 : std_logic_vector(0 to 0) := (others => '0');
    variable r7226 : std_logic_vector(0 to 0) := (others => '0');
    variable r7225 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r7226 := "1";
    null;
    r7227 := (r7226);
    r7228 := "1";
    null;
    r7229 := (r7228);
    r7230 := "0";
    null;
    r7231 := (r7230);
    r7232 := "0";
    null;
    r7233 := (r7232);
    r7234 := "0";
    null;
    r7235 := (r7234);
    r7236 := "1";
    null;
    r7237 := (r7236);
    r7238 := "1";
    null;
    r7239 := (r7238);
    r7240 := "0";
    null;
    r7241 := (r7240);
    r7242 := "0";
    null;
    r7243 := (r7242);
    r7244 := "1";
    null;
    r7245 := (r7244);
    r7246 := "1";
    null;
    r7247 := (r7246);
    r7248 := "1";
    null;
    r7249 := (r7248);
    r7250 := "0";
    null;
    r7251 := (r7250);
    r7252 := "0";
    null;
    r7253 := (r7252);
    r7254 := "0";
    null;
    r7255 := (r7254);
    r7256 := "1";
    null;
    r7257 := (r7256);
    r7258 := "0";
    null;
    r7259 := (r7258);
    r7260 := "1";
    null;
    r7261 := (r7260);
    r7262 := "1";
    null;
    r7263 := (r7262);
    r7264 := "1";
    null;
    r7265 := (r7264);
    r7266 := "1";
    null;
    r7267 := (r7266);
    r7268 := "0";
    null;
    r7269 := (r7268);
    r7270 := "0";
    null;
    r7271 := (r7270);
    r7272 := "0";
    null;
    r7273 := (r7272);
    r7274 := "1";
    null;
    r7275 := (r7274);
    r7276 := "1";
    null;
    r7277 := (r7276);
    r7278 := "1";
    null;
    r7279 := (r7278);
    r7280 := "1";
    null;
    r7281 := (r7280);
    r7282 := "0";
    null;
    r7283 := (r7282);
    r7284 := "0";
    null;
    r7285 := (r7284);
    r7286 := "1";
    null;
    r7287 := (r7286);
    r7288 := "0";
    null;
    r7289 := (r7288);
    r7225 := (r7227 & r7229 & r7231 & r7233 & r7235 & r7237 & r7239 & r7241 & r7243 & r7245 & r7247 & r7249 & r7251 & r7253 & r7255 & r7257 & r7259 & r7261 & r7263 & r7265 & r7267 & r7269 & r7271 & r7273 & r7275 & r7277 & r7279 & r7281 & r7283 & r7285 & r7287 & r7289);
    return r7225;
  end rewire_MetaprogrammingRWwc67178f2_7224;
  function rewire_MetaprogrammingRWwbef9a3f7_7155 return std_logic_vector
  is
    variable r7220 : std_logic_vector(0 to 0) := (others => '0');
    variable r7219 : std_logic_vector(0 to 0) := (others => '0');
    variable r7218 : std_logic_vector(0 to 0) := (others => '0');
    variable r7217 : std_logic_vector(0 to 0) := (others => '0');
    variable r7216 : std_logic_vector(0 to 0) := (others => '0');
    variable r7215 : std_logic_vector(0 to 0) := (others => '0');
    variable r7214 : std_logic_vector(0 to 0) := (others => '0');
    variable r7213 : std_logic_vector(0 to 0) := (others => '0');
    variable r7212 : std_logic_vector(0 to 0) := (others => '0');
    variable r7211 : std_logic_vector(0 to 0) := (others => '0');
    variable r7210 : std_logic_vector(0 to 0) := (others => '0');
    variable r7209 : std_logic_vector(0 to 0) := (others => '0');
    variable r7208 : std_logic_vector(0 to 0) := (others => '0');
    variable r7207 : std_logic_vector(0 to 0) := (others => '0');
    variable r7206 : std_logic_vector(0 to 0) := (others => '0');
    variable r7205 : std_logic_vector(0 to 0) := (others => '0');
    variable r7204 : std_logic_vector(0 to 0) := (others => '0');
    variable r7203 : std_logic_vector(0 to 0) := (others => '0');
    variable r7202 : std_logic_vector(0 to 0) := (others => '0');
    variable r7201 : std_logic_vector(0 to 0) := (others => '0');
    variable r7200 : std_logic_vector(0 to 0) := (others => '0');
    variable r7199 : std_logic_vector(0 to 0) := (others => '0');
    variable r7198 : std_logic_vector(0 to 0) := (others => '0');
    variable r7197 : std_logic_vector(0 to 0) := (others => '0');
    variable r7196 : std_logic_vector(0 to 0) := (others => '0');
    variable r7195 : std_logic_vector(0 to 0) := (others => '0');
    variable r7194 : std_logic_vector(0 to 0) := (others => '0');
    variable r7193 : std_logic_vector(0 to 0) := (others => '0');
    variable r7192 : std_logic_vector(0 to 0) := (others => '0');
    variable r7191 : std_logic_vector(0 to 0) := (others => '0');
    variable r7190 : std_logic_vector(0 to 0) := (others => '0');
    variable r7189 : std_logic_vector(0 to 0) := (others => '0');
    variable r7188 : std_logic_vector(0 to 0) := (others => '0');
    variable r7187 : std_logic_vector(0 to 0) := (others => '0');
    variable r7186 : std_logic_vector(0 to 0) := (others => '0');
    variable r7185 : std_logic_vector(0 to 0) := (others => '0');
    variable r7184 : std_logic_vector(0 to 0) := (others => '0');
    variable r7183 : std_logic_vector(0 to 0) := (others => '0');
    variable r7182 : std_logic_vector(0 to 0) := (others => '0');
    variable r7181 : std_logic_vector(0 to 0) := (others => '0');
    variable r7180 : std_logic_vector(0 to 0) := (others => '0');
    variable r7179 : std_logic_vector(0 to 0) := (others => '0');
    variable r7178 : std_logic_vector(0 to 0) := (others => '0');
    variable r7177 : std_logic_vector(0 to 0) := (others => '0');
    variable r7176 : std_logic_vector(0 to 0) := (others => '0');
    variable r7175 : std_logic_vector(0 to 0) := (others => '0');
    variable r7174 : std_logic_vector(0 to 0) := (others => '0');
    variable r7173 : std_logic_vector(0 to 0) := (others => '0');
    variable r7172 : std_logic_vector(0 to 0) := (others => '0');
    variable r7171 : std_logic_vector(0 to 0) := (others => '0');
    variable r7170 : std_logic_vector(0 to 0) := (others => '0');
    variable r7169 : std_logic_vector(0 to 0) := (others => '0');
    variable r7168 : std_logic_vector(0 to 0) := (others => '0');
    variable r7167 : std_logic_vector(0 to 0) := (others => '0');
    variable r7166 : std_logic_vector(0 to 0) := (others => '0');
    variable r7165 : std_logic_vector(0 to 0) := (others => '0');
    variable r7164 : std_logic_vector(0 to 0) := (others => '0');
    variable r7163 : std_logic_vector(0 to 0) := (others => '0');
    variable r7162 : std_logic_vector(0 to 0) := (others => '0');
    variable r7161 : std_logic_vector(0 to 0) := (others => '0');
    variable r7160 : std_logic_vector(0 to 0) := (others => '0');
    variable r7159 : std_logic_vector(0 to 0) := (others => '0');
    variable r7158 : std_logic_vector(0 to 0) := (others => '0');
    variable r7157 : std_logic_vector(0 to 0) := (others => '0');
    variable r7156 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r7157 := "1";
    null;
    r7158 := (r7157);
    r7159 := "0";
    null;
    r7160 := (r7159);
    r7161 := "1";
    null;
    r7162 := (r7161);
    r7163 := "1";
    null;
    r7164 := (r7163);
    r7165 := "1";
    null;
    r7166 := (r7165);
    r7167 := "1";
    null;
    r7168 := (r7167);
    r7169 := "1";
    null;
    r7170 := (r7169);
    r7171 := "0";
    null;
    r7172 := (r7171);
    r7173 := "1";
    null;
    r7174 := (r7173);
    r7175 := "1";
    null;
    r7176 := (r7175);
    r7177 := "1";
    null;
    r7178 := (r7177);
    r7179 := "1";
    null;
    r7180 := (r7179);
    r7181 := "1";
    null;
    r7182 := (r7181);
    r7183 := "0";
    null;
    r7184 := (r7183);
    r7185 := "0";
    null;
    r7186 := (r7185);
    r7187 := "1";
    null;
    r7188 := (r7187);
    r7189 := "1";
    null;
    r7190 := (r7189);
    r7191 := "0";
    null;
    r7192 := (r7191);
    r7193 := "1";
    null;
    r7194 := (r7193);
    r7195 := "0";
    null;
    r7196 := (r7195);
    r7197 := "0";
    null;
    r7198 := (r7197);
    r7199 := "0";
    null;
    r7200 := (r7199);
    r7201 := "1";
    null;
    r7202 := (r7201);
    r7203 := "1";
    null;
    r7204 := (r7203);
    r7205 := "1";
    null;
    r7206 := (r7205);
    r7207 := "1";
    null;
    r7208 := (r7207);
    r7209 := "1";
    null;
    r7210 := (r7209);
    r7211 := "1";
    null;
    r7212 := (r7211);
    r7213 := "0";
    null;
    r7214 := (r7213);
    r7215 := "1";
    null;
    r7216 := (r7215);
    r7217 := "1";
    null;
    r7218 := (r7217);
    r7219 := "1";
    null;
    r7220 := (r7219);
    r7156 := (r7158 & r7160 & r7162 & r7164 & r7166 & r7168 & r7170 & r7172 & r7174 & r7176 & r7178 & r7180 & r7182 & r7184 & r7186 & r7188 & r7190 & r7192 & r7194 & r7196 & r7198 & r7200 & r7202 & r7204 & r7206 & r7208 & r7210 & r7212 & r7214 & r7216 & r7218 & r7220);
    return r7156;
  end rewire_MetaprogrammingRWwbef9a3f7_7155;
  function rewire_MetaprogrammingRWwa4506ceb_7086 return std_logic_vector
  is
    variable r7151 : std_logic_vector(0 to 0) := (others => '0');
    variable r7150 : std_logic_vector(0 to 0) := (others => '0');
    variable r7149 : std_logic_vector(0 to 0) := (others => '0');
    variable r7148 : std_logic_vector(0 to 0) := (others => '0');
    variable r7147 : std_logic_vector(0 to 0) := (others => '0');
    variable r7146 : std_logic_vector(0 to 0) := (others => '0');
    variable r7145 : std_logic_vector(0 to 0) := (others => '0');
    variable r7144 : std_logic_vector(0 to 0) := (others => '0');
    variable r7143 : std_logic_vector(0 to 0) := (others => '0');
    variable r7142 : std_logic_vector(0 to 0) := (others => '0');
    variable r7141 : std_logic_vector(0 to 0) := (others => '0');
    variable r7140 : std_logic_vector(0 to 0) := (others => '0');
    variable r7139 : std_logic_vector(0 to 0) := (others => '0');
    variable r7138 : std_logic_vector(0 to 0) := (others => '0');
    variable r7137 : std_logic_vector(0 to 0) := (others => '0');
    variable r7136 : std_logic_vector(0 to 0) := (others => '0');
    variable r7135 : std_logic_vector(0 to 0) := (others => '0');
    variable r7134 : std_logic_vector(0 to 0) := (others => '0');
    variable r7133 : std_logic_vector(0 to 0) := (others => '0');
    variable r7132 : std_logic_vector(0 to 0) := (others => '0');
    variable r7131 : std_logic_vector(0 to 0) := (others => '0');
    variable r7130 : std_logic_vector(0 to 0) := (others => '0');
    variable r7129 : std_logic_vector(0 to 0) := (others => '0');
    variable r7128 : std_logic_vector(0 to 0) := (others => '0');
    variable r7127 : std_logic_vector(0 to 0) := (others => '0');
    variable r7126 : std_logic_vector(0 to 0) := (others => '0');
    variable r7125 : std_logic_vector(0 to 0) := (others => '0');
    variable r7124 : std_logic_vector(0 to 0) := (others => '0');
    variable r7123 : std_logic_vector(0 to 0) := (others => '0');
    variable r7122 : std_logic_vector(0 to 0) := (others => '0');
    variable r7121 : std_logic_vector(0 to 0) := (others => '0');
    variable r7120 : std_logic_vector(0 to 0) := (others => '0');
    variable r7119 : std_logic_vector(0 to 0) := (others => '0');
    variable r7118 : std_logic_vector(0 to 0) := (others => '0');
    variable r7117 : std_logic_vector(0 to 0) := (others => '0');
    variable r7116 : std_logic_vector(0 to 0) := (others => '0');
    variable r7115 : std_logic_vector(0 to 0) := (others => '0');
    variable r7114 : std_logic_vector(0 to 0) := (others => '0');
    variable r7113 : std_logic_vector(0 to 0) := (others => '0');
    variable r7112 : std_logic_vector(0 to 0) := (others => '0');
    variable r7111 : std_logic_vector(0 to 0) := (others => '0');
    variable r7110 : std_logic_vector(0 to 0) := (others => '0');
    variable r7109 : std_logic_vector(0 to 0) := (others => '0');
    variable r7108 : std_logic_vector(0 to 0) := (others => '0');
    variable r7107 : std_logic_vector(0 to 0) := (others => '0');
    variable r7106 : std_logic_vector(0 to 0) := (others => '0');
    variable r7105 : std_logic_vector(0 to 0) := (others => '0');
    variable r7104 : std_logic_vector(0 to 0) := (others => '0');
    variable r7103 : std_logic_vector(0 to 0) := (others => '0');
    variable r7102 : std_logic_vector(0 to 0) := (others => '0');
    variable r7101 : std_logic_vector(0 to 0) := (others => '0');
    variable r7100 : std_logic_vector(0 to 0) := (others => '0');
    variable r7099 : std_logic_vector(0 to 0) := (others => '0');
    variable r7098 : std_logic_vector(0 to 0) := (others => '0');
    variable r7097 : std_logic_vector(0 to 0) := (others => '0');
    variable r7096 : std_logic_vector(0 to 0) := (others => '0');
    variable r7095 : std_logic_vector(0 to 0) := (others => '0');
    variable r7094 : std_logic_vector(0 to 0) := (others => '0');
    variable r7093 : std_logic_vector(0 to 0) := (others => '0');
    variable r7092 : std_logic_vector(0 to 0) := (others => '0');
    variable r7091 : std_logic_vector(0 to 0) := (others => '0');
    variable r7090 : std_logic_vector(0 to 0) := (others => '0');
    variable r7089 : std_logic_vector(0 to 0) := (others => '0');
    variable r7088 : std_logic_vector(0 to 0) := (others => '0');
    variable r7087 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r7088 := "1";
    null;
    r7089 := (r7088);
    r7090 := "0";
    null;
    r7091 := (r7090);
    r7092 := "1";
    null;
    r7093 := (r7092);
    r7094 := "0";
    null;
    r7095 := (r7094);
    r7096 := "0";
    null;
    r7097 := (r7096);
    r7098 := "1";
    null;
    r7099 := (r7098);
    r7100 := "0";
    null;
    r7101 := (r7100);
    r7102 := "0";
    null;
    r7103 := (r7102);
    r7104 := "0";
    null;
    r7105 := (r7104);
    r7106 := "1";
    null;
    r7107 := (r7106);
    r7108 := "0";
    null;
    r7109 := (r7108);
    r7110 := "1";
    null;
    r7111 := (r7110);
    r7112 := "0";
    null;
    r7113 := (r7112);
    r7114 := "0";
    null;
    r7115 := (r7114);
    r7116 := "0";
    null;
    r7117 := (r7116);
    r7118 := "0";
    null;
    r7119 := (r7118);
    r7120 := "0";
    null;
    r7121 := (r7120);
    r7122 := "1";
    null;
    r7123 := (r7122);
    r7124 := "1";
    null;
    r7125 := (r7124);
    r7126 := "0";
    null;
    r7127 := (r7126);
    r7128 := "1";
    null;
    r7129 := (r7128);
    r7130 := "1";
    null;
    r7131 := (r7130);
    r7132 := "0";
    null;
    r7133 := (r7132);
    r7134 := "0";
    null;
    r7135 := (r7134);
    r7136 := "1";
    null;
    r7137 := (r7136);
    r7138 := "1";
    null;
    r7139 := (r7138);
    r7140 := "1";
    null;
    r7141 := (r7140);
    r7142 := "0";
    null;
    r7143 := (r7142);
    r7144 := "1";
    null;
    r7145 := (r7144);
    r7146 := "0";
    null;
    r7147 := (r7146);
    r7148 := "1";
    null;
    r7149 := (r7148);
    r7150 := "1";
    null;
    r7151 := (r7150);
    r7087 := (r7089 & r7091 & r7093 & r7095 & r7097 & r7099 & r7101 & r7103 & r7105 & r7107 & r7109 & r7111 & r7113 & r7115 & r7117 & r7119 & r7121 & r7123 & r7125 & r7127 & r7129 & r7131 & r7133 & r7135 & r7137 & r7139 & r7141 & r7143 & r7145 & r7147 & r7149 & r7151);
    return r7087;
  end rewire_MetaprogrammingRWwa4506ceb_7086;
  function rewire_MetaprogrammingRWw90befffa_7017 return std_logic_vector
  is
    variable r7082 : std_logic_vector(0 to 0) := (others => '0');
    variable r7081 : std_logic_vector(0 to 0) := (others => '0');
    variable r7080 : std_logic_vector(0 to 0) := (others => '0');
    variable r7079 : std_logic_vector(0 to 0) := (others => '0');
    variable r7078 : std_logic_vector(0 to 0) := (others => '0');
    variable r7077 : std_logic_vector(0 to 0) := (others => '0');
    variable r7076 : std_logic_vector(0 to 0) := (others => '0');
    variable r7075 : std_logic_vector(0 to 0) := (others => '0');
    variable r7074 : std_logic_vector(0 to 0) := (others => '0');
    variable r7073 : std_logic_vector(0 to 0) := (others => '0');
    variable r7072 : std_logic_vector(0 to 0) := (others => '0');
    variable r7071 : std_logic_vector(0 to 0) := (others => '0');
    variable r7070 : std_logic_vector(0 to 0) := (others => '0');
    variable r7069 : std_logic_vector(0 to 0) := (others => '0');
    variable r7068 : std_logic_vector(0 to 0) := (others => '0');
    variable r7067 : std_logic_vector(0 to 0) := (others => '0');
    variable r7066 : std_logic_vector(0 to 0) := (others => '0');
    variable r7065 : std_logic_vector(0 to 0) := (others => '0');
    variable r7064 : std_logic_vector(0 to 0) := (others => '0');
    variable r7063 : std_logic_vector(0 to 0) := (others => '0');
    variable r7062 : std_logic_vector(0 to 0) := (others => '0');
    variable r7061 : std_logic_vector(0 to 0) := (others => '0');
    variable r7060 : std_logic_vector(0 to 0) := (others => '0');
    variable r7059 : std_logic_vector(0 to 0) := (others => '0');
    variable r7058 : std_logic_vector(0 to 0) := (others => '0');
    variable r7057 : std_logic_vector(0 to 0) := (others => '0');
    variable r7056 : std_logic_vector(0 to 0) := (others => '0');
    variable r7055 : std_logic_vector(0 to 0) := (others => '0');
    variable r7054 : std_logic_vector(0 to 0) := (others => '0');
    variable r7053 : std_logic_vector(0 to 0) := (others => '0');
    variable r7052 : std_logic_vector(0 to 0) := (others => '0');
    variable r7051 : std_logic_vector(0 to 0) := (others => '0');
    variable r7050 : std_logic_vector(0 to 0) := (others => '0');
    variable r7049 : std_logic_vector(0 to 0) := (others => '0');
    variable r7048 : std_logic_vector(0 to 0) := (others => '0');
    variable r7047 : std_logic_vector(0 to 0) := (others => '0');
    variable r7046 : std_logic_vector(0 to 0) := (others => '0');
    variable r7045 : std_logic_vector(0 to 0) := (others => '0');
    variable r7044 : std_logic_vector(0 to 0) := (others => '0');
    variable r7043 : std_logic_vector(0 to 0) := (others => '0');
    variable r7042 : std_logic_vector(0 to 0) := (others => '0');
    variable r7041 : std_logic_vector(0 to 0) := (others => '0');
    variable r7040 : std_logic_vector(0 to 0) := (others => '0');
    variable r7039 : std_logic_vector(0 to 0) := (others => '0');
    variable r7038 : std_logic_vector(0 to 0) := (others => '0');
    variable r7037 : std_logic_vector(0 to 0) := (others => '0');
    variable r7036 : std_logic_vector(0 to 0) := (others => '0');
    variable r7035 : std_logic_vector(0 to 0) := (others => '0');
    variable r7034 : std_logic_vector(0 to 0) := (others => '0');
    variable r7033 : std_logic_vector(0 to 0) := (others => '0');
    variable r7032 : std_logic_vector(0 to 0) := (others => '0');
    variable r7031 : std_logic_vector(0 to 0) := (others => '0');
    variable r7030 : std_logic_vector(0 to 0) := (others => '0');
    variable r7029 : std_logic_vector(0 to 0) := (others => '0');
    variable r7028 : std_logic_vector(0 to 0) := (others => '0');
    variable r7027 : std_logic_vector(0 to 0) := (others => '0');
    variable r7026 : std_logic_vector(0 to 0) := (others => '0');
    variable r7025 : std_logic_vector(0 to 0) := (others => '0');
    variable r7024 : std_logic_vector(0 to 0) := (others => '0');
    variable r7023 : std_logic_vector(0 to 0) := (others => '0');
    variable r7022 : std_logic_vector(0 to 0) := (others => '0');
    variable r7021 : std_logic_vector(0 to 0) := (others => '0');
    variable r7020 : std_logic_vector(0 to 0) := (others => '0');
    variable r7019 : std_logic_vector(0 to 0) := (others => '0');
    variable r7018 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r7019 := "1";
    null;
    r7020 := (r7019);
    r7021 := "0";
    null;
    r7022 := (r7021);
    r7023 := "0";
    null;
    r7024 := (r7023);
    r7025 := "1";
    null;
    r7026 := (r7025);
    r7027 := "0";
    null;
    r7028 := (r7027);
    r7029 := "0";
    null;
    r7030 := (r7029);
    r7031 := "0";
    null;
    r7032 := (r7031);
    r7033 := "0";
    null;
    r7034 := (r7033);
    r7035 := "1";
    null;
    r7036 := (r7035);
    r7037 := "0";
    null;
    r7038 := (r7037);
    r7039 := "1";
    null;
    r7040 := (r7039);
    r7041 := "1";
    null;
    r7042 := (r7041);
    r7043 := "1";
    null;
    r7044 := (r7043);
    r7045 := "1";
    null;
    r7046 := (r7045);
    r7047 := "1";
    null;
    r7048 := (r7047);
    r7049 := "0";
    null;
    r7050 := (r7049);
    r7051 := "1";
    null;
    r7052 := (r7051);
    r7053 := "1";
    null;
    r7054 := (r7053);
    r7055 := "1";
    null;
    r7056 := (r7055);
    r7057 := "1";
    null;
    r7058 := (r7057);
    r7059 := "1";
    null;
    r7060 := (r7059);
    r7061 := "1";
    null;
    r7062 := (r7061);
    r7063 := "1";
    null;
    r7064 := (r7063);
    r7065 := "1";
    null;
    r7066 := (r7065);
    r7067 := "1";
    null;
    r7068 := (r7067);
    r7069 := "1";
    null;
    r7070 := (r7069);
    r7071 := "1";
    null;
    r7072 := (r7071);
    r7073 := "1";
    null;
    r7074 := (r7073);
    r7075 := "1";
    null;
    r7076 := (r7075);
    r7077 := "0";
    null;
    r7078 := (r7077);
    r7079 := "1";
    null;
    r7080 := (r7079);
    r7081 := "0";
    null;
    r7082 := (r7081);
    r7018 := (r7020 & r7022 & r7024 & r7026 & r7028 & r7030 & r7032 & r7034 & r7036 & r7038 & r7040 & r7042 & r7044 & r7046 & r7048 & r7050 & r7052 & r7054 & r7056 & r7058 & r7060 & r7062 & r7064 & r7066 & r7068 & r7070 & r7072 & r7074 & r7076 & r7078 & r7080 & r7082);
    return r7018;
  end rewire_MetaprogrammingRWw90befffa_7017;
  function rewire_MetaprogrammingRWw8cc70208_6948 return std_logic_vector
  is
    variable r7013 : std_logic_vector(0 to 0) := (others => '0');
    variable r7012 : std_logic_vector(0 to 0) := (others => '0');
    variable r7011 : std_logic_vector(0 to 0) := (others => '0');
    variable r7010 : std_logic_vector(0 to 0) := (others => '0');
    variable r7009 : std_logic_vector(0 to 0) := (others => '0');
    variable r7008 : std_logic_vector(0 to 0) := (others => '0');
    variable r7007 : std_logic_vector(0 to 0) := (others => '0');
    variable r7006 : std_logic_vector(0 to 0) := (others => '0');
    variable r7005 : std_logic_vector(0 to 0) := (others => '0');
    variable r7004 : std_logic_vector(0 to 0) := (others => '0');
    variable r7003 : std_logic_vector(0 to 0) := (others => '0');
    variable r7002 : std_logic_vector(0 to 0) := (others => '0');
    variable r7001 : std_logic_vector(0 to 0) := (others => '0');
    variable r7000 : std_logic_vector(0 to 0) := (others => '0');
    variable r6999 : std_logic_vector(0 to 0) := (others => '0');
    variable r6998 : std_logic_vector(0 to 0) := (others => '0');
    variable r6997 : std_logic_vector(0 to 0) := (others => '0');
    variable r6996 : std_logic_vector(0 to 0) := (others => '0');
    variable r6995 : std_logic_vector(0 to 0) := (others => '0');
    variable r6994 : std_logic_vector(0 to 0) := (others => '0');
    variable r6993 : std_logic_vector(0 to 0) := (others => '0');
    variable r6992 : std_logic_vector(0 to 0) := (others => '0');
    variable r6991 : std_logic_vector(0 to 0) := (others => '0');
    variable r6990 : std_logic_vector(0 to 0) := (others => '0');
    variable r6989 : std_logic_vector(0 to 0) := (others => '0');
    variable r6988 : std_logic_vector(0 to 0) := (others => '0');
    variable r6987 : std_logic_vector(0 to 0) := (others => '0');
    variable r6986 : std_logic_vector(0 to 0) := (others => '0');
    variable r6985 : std_logic_vector(0 to 0) := (others => '0');
    variable r6984 : std_logic_vector(0 to 0) := (others => '0');
    variable r6983 : std_logic_vector(0 to 0) := (others => '0');
    variable r6982 : std_logic_vector(0 to 0) := (others => '0');
    variable r6981 : std_logic_vector(0 to 0) := (others => '0');
    variable r6980 : std_logic_vector(0 to 0) := (others => '0');
    variable r6979 : std_logic_vector(0 to 0) := (others => '0');
    variable r6978 : std_logic_vector(0 to 0) := (others => '0');
    variable r6977 : std_logic_vector(0 to 0) := (others => '0');
    variable r6976 : std_logic_vector(0 to 0) := (others => '0');
    variable r6975 : std_logic_vector(0 to 0) := (others => '0');
    variable r6974 : std_logic_vector(0 to 0) := (others => '0');
    variable r6973 : std_logic_vector(0 to 0) := (others => '0');
    variable r6972 : std_logic_vector(0 to 0) := (others => '0');
    variable r6971 : std_logic_vector(0 to 0) := (others => '0');
    variable r6970 : std_logic_vector(0 to 0) := (others => '0');
    variable r6969 : std_logic_vector(0 to 0) := (others => '0');
    variable r6968 : std_logic_vector(0 to 0) := (others => '0');
    variable r6967 : std_logic_vector(0 to 0) := (others => '0');
    variable r6966 : std_logic_vector(0 to 0) := (others => '0');
    variable r6965 : std_logic_vector(0 to 0) := (others => '0');
    variable r6964 : std_logic_vector(0 to 0) := (others => '0');
    variable r6963 : std_logic_vector(0 to 0) := (others => '0');
    variable r6962 : std_logic_vector(0 to 0) := (others => '0');
    variable r6961 : std_logic_vector(0 to 0) := (others => '0');
    variable r6960 : std_logic_vector(0 to 0) := (others => '0');
    variable r6959 : std_logic_vector(0 to 0) := (others => '0');
    variable r6958 : std_logic_vector(0 to 0) := (others => '0');
    variable r6957 : std_logic_vector(0 to 0) := (others => '0');
    variable r6956 : std_logic_vector(0 to 0) := (others => '0');
    variable r6955 : std_logic_vector(0 to 0) := (others => '0');
    variable r6954 : std_logic_vector(0 to 0) := (others => '0');
    variable r6953 : std_logic_vector(0 to 0) := (others => '0');
    variable r6952 : std_logic_vector(0 to 0) := (others => '0');
    variable r6951 : std_logic_vector(0 to 0) := (others => '0');
    variable r6950 : std_logic_vector(0 to 0) := (others => '0');
    variable r6949 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r6950 := "1";
    null;
    r6951 := (r6950);
    r6952 := "0";
    null;
    r6953 := (r6952);
    r6954 := "0";
    null;
    r6955 := (r6954);
    r6956 := "0";
    null;
    r6957 := (r6956);
    r6958 := "1";
    null;
    r6959 := (r6958);
    r6960 := "1";
    null;
    r6961 := (r6960);
    r6962 := "0";
    null;
    r6963 := (r6962);
    r6964 := "0";
    null;
    r6965 := (r6964);
    r6966 := "1";
    null;
    r6967 := (r6966);
    r6968 := "1";
    null;
    r6969 := (r6968);
    r6970 := "0";
    null;
    r6971 := (r6970);
    r6972 := "0";
    null;
    r6973 := (r6972);
    r6974 := "0";
    null;
    r6975 := (r6974);
    r6976 := "1";
    null;
    r6977 := (r6976);
    r6978 := "1";
    null;
    r6979 := (r6978);
    r6980 := "1";
    null;
    r6981 := (r6980);
    r6982 := "0";
    null;
    r6983 := (r6982);
    r6984 := "0";
    null;
    r6985 := (r6984);
    r6986 := "0";
    null;
    r6987 := (r6986);
    r6988 := "0";
    null;
    r6989 := (r6988);
    r6990 := "0";
    null;
    r6991 := (r6990);
    r6992 := "0";
    null;
    r6993 := (r6992);
    r6994 := "1";
    null;
    r6995 := (r6994);
    r6996 := "0";
    null;
    r6997 := (r6996);
    r6998 := "0";
    null;
    r6999 := (r6998);
    r7000 := "0";
    null;
    r7001 := (r7000);
    r7002 := "0";
    null;
    r7003 := (r7002);
    r7004 := "0";
    null;
    r7005 := (r7004);
    r7006 := "1";
    null;
    r7007 := (r7006);
    r7008 := "0";
    null;
    r7009 := (r7008);
    r7010 := "0";
    null;
    r7011 := (r7010);
    r7012 := "0";
    null;
    r7013 := (r7012);
    r6949 := (r6951 & r6953 & r6955 & r6957 & r6959 & r6961 & r6963 & r6965 & r6967 & r6969 & r6971 & r6973 & r6975 & r6977 & r6979 & r6981 & r6983 & r6985 & r6987 & r6989 & r6991 & r6993 & r6995 & r6997 & r6999 & r7001 & r7003 & r7005 & r7007 & r7009 & r7011 & r7013);
    return r6949;
  end rewire_MetaprogrammingRWw8cc70208_6948;
  function rewire_MetaprogrammingRWw84c87814_6879 return std_logic_vector
  is
    variable r6944 : std_logic_vector(0 to 0) := (others => '0');
    variable r6943 : std_logic_vector(0 to 0) := (others => '0');
    variable r6942 : std_logic_vector(0 to 0) := (others => '0');
    variable r6941 : std_logic_vector(0 to 0) := (others => '0');
    variable r6940 : std_logic_vector(0 to 0) := (others => '0');
    variable r6939 : std_logic_vector(0 to 0) := (others => '0');
    variable r6938 : std_logic_vector(0 to 0) := (others => '0');
    variable r6937 : std_logic_vector(0 to 0) := (others => '0');
    variable r6936 : std_logic_vector(0 to 0) := (others => '0');
    variable r6935 : std_logic_vector(0 to 0) := (others => '0');
    variable r6934 : std_logic_vector(0 to 0) := (others => '0');
    variable r6933 : std_logic_vector(0 to 0) := (others => '0');
    variable r6932 : std_logic_vector(0 to 0) := (others => '0');
    variable r6931 : std_logic_vector(0 to 0) := (others => '0');
    variable r6930 : std_logic_vector(0 to 0) := (others => '0');
    variable r6929 : std_logic_vector(0 to 0) := (others => '0');
    variable r6928 : std_logic_vector(0 to 0) := (others => '0');
    variable r6927 : std_logic_vector(0 to 0) := (others => '0');
    variable r6926 : std_logic_vector(0 to 0) := (others => '0');
    variable r6925 : std_logic_vector(0 to 0) := (others => '0');
    variable r6924 : std_logic_vector(0 to 0) := (others => '0');
    variable r6923 : std_logic_vector(0 to 0) := (others => '0');
    variable r6922 : std_logic_vector(0 to 0) := (others => '0');
    variable r6921 : std_logic_vector(0 to 0) := (others => '0');
    variable r6920 : std_logic_vector(0 to 0) := (others => '0');
    variable r6919 : std_logic_vector(0 to 0) := (others => '0');
    variable r6918 : std_logic_vector(0 to 0) := (others => '0');
    variable r6917 : std_logic_vector(0 to 0) := (others => '0');
    variable r6916 : std_logic_vector(0 to 0) := (others => '0');
    variable r6915 : std_logic_vector(0 to 0) := (others => '0');
    variable r6914 : std_logic_vector(0 to 0) := (others => '0');
    variable r6913 : std_logic_vector(0 to 0) := (others => '0');
    variable r6912 : std_logic_vector(0 to 0) := (others => '0');
    variable r6911 : std_logic_vector(0 to 0) := (others => '0');
    variable r6910 : std_logic_vector(0 to 0) := (others => '0');
    variable r6909 : std_logic_vector(0 to 0) := (others => '0');
    variable r6908 : std_logic_vector(0 to 0) := (others => '0');
    variable r6907 : std_logic_vector(0 to 0) := (others => '0');
    variable r6906 : std_logic_vector(0 to 0) := (others => '0');
    variable r6905 : std_logic_vector(0 to 0) := (others => '0');
    variable r6904 : std_logic_vector(0 to 0) := (others => '0');
    variable r6903 : std_logic_vector(0 to 0) := (others => '0');
    variable r6902 : std_logic_vector(0 to 0) := (others => '0');
    variable r6901 : std_logic_vector(0 to 0) := (others => '0');
    variable r6900 : std_logic_vector(0 to 0) := (others => '0');
    variable r6899 : std_logic_vector(0 to 0) := (others => '0');
    variable r6898 : std_logic_vector(0 to 0) := (others => '0');
    variable r6897 : std_logic_vector(0 to 0) := (others => '0');
    variable r6896 : std_logic_vector(0 to 0) := (others => '0');
    variable r6895 : std_logic_vector(0 to 0) := (others => '0');
    variable r6894 : std_logic_vector(0 to 0) := (others => '0');
    variable r6893 : std_logic_vector(0 to 0) := (others => '0');
    variable r6892 : std_logic_vector(0 to 0) := (others => '0');
    variable r6891 : std_logic_vector(0 to 0) := (others => '0');
    variable r6890 : std_logic_vector(0 to 0) := (others => '0');
    variable r6889 : std_logic_vector(0 to 0) := (others => '0');
    variable r6888 : std_logic_vector(0 to 0) := (others => '0');
    variable r6887 : std_logic_vector(0 to 0) := (others => '0');
    variable r6886 : std_logic_vector(0 to 0) := (others => '0');
    variable r6885 : std_logic_vector(0 to 0) := (others => '0');
    variable r6884 : std_logic_vector(0 to 0) := (others => '0');
    variable r6883 : std_logic_vector(0 to 0) := (others => '0');
    variable r6882 : std_logic_vector(0 to 0) := (others => '0');
    variable r6881 : std_logic_vector(0 to 0) := (others => '0');
    variable r6880 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r6881 := "1";
    null;
    r6882 := (r6881);
    r6883 := "0";
    null;
    r6884 := (r6883);
    r6885 := "0";
    null;
    r6886 := (r6885);
    r6887 := "0";
    null;
    r6888 := (r6887);
    r6889 := "0";
    null;
    r6890 := (r6889);
    r6891 := "1";
    null;
    r6892 := (r6891);
    r6893 := "0";
    null;
    r6894 := (r6893);
    r6895 := "0";
    null;
    r6896 := (r6895);
    r6897 := "1";
    null;
    r6898 := (r6897);
    r6899 := "1";
    null;
    r6900 := (r6899);
    r6901 := "0";
    null;
    r6902 := (r6901);
    r6903 := "0";
    null;
    r6904 := (r6903);
    r6905 := "1";
    null;
    r6906 := (r6905);
    r6907 := "0";
    null;
    r6908 := (r6907);
    r6909 := "0";
    null;
    r6910 := (r6909);
    r6911 := "0";
    null;
    r6912 := (r6911);
    r6913 := "0";
    null;
    r6914 := (r6913);
    r6915 := "1";
    null;
    r6916 := (r6915);
    r6917 := "1";
    null;
    r6918 := (r6917);
    r6919 := "1";
    null;
    r6920 := (r6919);
    r6921 := "1";
    null;
    r6922 := (r6921);
    r6923 := "0";
    null;
    r6924 := (r6923);
    r6925 := "0";
    null;
    r6926 := (r6925);
    r6927 := "0";
    null;
    r6928 := (r6927);
    r6929 := "0";
    null;
    r6930 := (r6929);
    r6931 := "0";
    null;
    r6932 := (r6931);
    r6933 := "0";
    null;
    r6934 := (r6933);
    r6935 := "1";
    null;
    r6936 := (r6935);
    r6937 := "0";
    null;
    r6938 := (r6937);
    r6939 := "1";
    null;
    r6940 := (r6939);
    r6941 := "0";
    null;
    r6942 := (r6941);
    r6943 := "0";
    null;
    r6944 := (r6943);
    r6880 := (r6882 & r6884 & r6886 & r6888 & r6890 & r6892 & r6894 & r6896 & r6898 & r6900 & r6902 & r6904 & r6906 & r6908 & r6910 & r6912 & r6914 & r6916 & r6918 & r6920 & r6922 & r6924 & r6926 & r6928 & r6930 & r6932 & r6934 & r6936 & r6938 & r6940 & r6942 & r6944);
    return r6880;
  end rewire_MetaprogrammingRWw84c87814_6879;
  function rewire_MetaprogrammingRWw78a5636f_6810 return std_logic_vector
  is
    variable r6875 : std_logic_vector(0 to 0) := (others => '0');
    variable r6874 : std_logic_vector(0 to 0) := (others => '0');
    variable r6873 : std_logic_vector(0 to 0) := (others => '0');
    variable r6872 : std_logic_vector(0 to 0) := (others => '0');
    variable r6871 : std_logic_vector(0 to 0) := (others => '0');
    variable r6870 : std_logic_vector(0 to 0) := (others => '0');
    variable r6869 : std_logic_vector(0 to 0) := (others => '0');
    variable r6868 : std_logic_vector(0 to 0) := (others => '0');
    variable r6867 : std_logic_vector(0 to 0) := (others => '0');
    variable r6866 : std_logic_vector(0 to 0) := (others => '0');
    variable r6865 : std_logic_vector(0 to 0) := (others => '0');
    variable r6864 : std_logic_vector(0 to 0) := (others => '0');
    variable r6863 : std_logic_vector(0 to 0) := (others => '0');
    variable r6862 : std_logic_vector(0 to 0) := (others => '0');
    variable r6861 : std_logic_vector(0 to 0) := (others => '0');
    variable r6860 : std_logic_vector(0 to 0) := (others => '0');
    variable r6859 : std_logic_vector(0 to 0) := (others => '0');
    variable r6858 : std_logic_vector(0 to 0) := (others => '0');
    variable r6857 : std_logic_vector(0 to 0) := (others => '0');
    variable r6856 : std_logic_vector(0 to 0) := (others => '0');
    variable r6855 : std_logic_vector(0 to 0) := (others => '0');
    variable r6854 : std_logic_vector(0 to 0) := (others => '0');
    variable r6853 : std_logic_vector(0 to 0) := (others => '0');
    variable r6852 : std_logic_vector(0 to 0) := (others => '0');
    variable r6851 : std_logic_vector(0 to 0) := (others => '0');
    variable r6850 : std_logic_vector(0 to 0) := (others => '0');
    variable r6849 : std_logic_vector(0 to 0) := (others => '0');
    variable r6848 : std_logic_vector(0 to 0) := (others => '0');
    variable r6847 : std_logic_vector(0 to 0) := (others => '0');
    variable r6846 : std_logic_vector(0 to 0) := (others => '0');
    variable r6845 : std_logic_vector(0 to 0) := (others => '0');
    variable r6844 : std_logic_vector(0 to 0) := (others => '0');
    variable r6843 : std_logic_vector(0 to 0) := (others => '0');
    variable r6842 : std_logic_vector(0 to 0) := (others => '0');
    variable r6841 : std_logic_vector(0 to 0) := (others => '0');
    variable r6840 : std_logic_vector(0 to 0) := (others => '0');
    variable r6839 : std_logic_vector(0 to 0) := (others => '0');
    variable r6838 : std_logic_vector(0 to 0) := (others => '0');
    variable r6837 : std_logic_vector(0 to 0) := (others => '0');
    variable r6836 : std_logic_vector(0 to 0) := (others => '0');
    variable r6835 : std_logic_vector(0 to 0) := (others => '0');
    variable r6834 : std_logic_vector(0 to 0) := (others => '0');
    variable r6833 : std_logic_vector(0 to 0) := (others => '0');
    variable r6832 : std_logic_vector(0 to 0) := (others => '0');
    variable r6831 : std_logic_vector(0 to 0) := (others => '0');
    variable r6830 : std_logic_vector(0 to 0) := (others => '0');
    variable r6829 : std_logic_vector(0 to 0) := (others => '0');
    variable r6828 : std_logic_vector(0 to 0) := (others => '0');
    variable r6827 : std_logic_vector(0 to 0) := (others => '0');
    variable r6826 : std_logic_vector(0 to 0) := (others => '0');
    variable r6825 : std_logic_vector(0 to 0) := (others => '0');
    variable r6824 : std_logic_vector(0 to 0) := (others => '0');
    variable r6823 : std_logic_vector(0 to 0) := (others => '0');
    variable r6822 : std_logic_vector(0 to 0) := (others => '0');
    variable r6821 : std_logic_vector(0 to 0) := (others => '0');
    variable r6820 : std_logic_vector(0 to 0) := (others => '0');
    variable r6819 : std_logic_vector(0 to 0) := (others => '0');
    variable r6818 : std_logic_vector(0 to 0) := (others => '0');
    variable r6817 : std_logic_vector(0 to 0) := (others => '0');
    variable r6816 : std_logic_vector(0 to 0) := (others => '0');
    variable r6815 : std_logic_vector(0 to 0) := (others => '0');
    variable r6814 : std_logic_vector(0 to 0) := (others => '0');
    variable r6813 : std_logic_vector(0 to 0) := (others => '0');
    variable r6812 : std_logic_vector(0 to 0) := (others => '0');
    variable r6811 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r6812 := "0";
    null;
    r6813 := (r6812);
    r6814 := "1";
    null;
    r6815 := (r6814);
    r6816 := "1";
    null;
    r6817 := (r6816);
    r6818 := "1";
    null;
    r6819 := (r6818);
    r6820 := "1";
    null;
    r6821 := (r6820);
    r6822 := "0";
    null;
    r6823 := (r6822);
    r6824 := "0";
    null;
    r6825 := (r6824);
    r6826 := "0";
    null;
    r6827 := (r6826);
    r6828 := "1";
    null;
    r6829 := (r6828);
    r6830 := "0";
    null;
    r6831 := (r6830);
    r6832 := "1";
    null;
    r6833 := (r6832);
    r6834 := "0";
    null;
    r6835 := (r6834);
    r6836 := "0";
    null;
    r6837 := (r6836);
    r6838 := "1";
    null;
    r6839 := (r6838);
    r6840 := "0";
    null;
    r6841 := (r6840);
    r6842 := "1";
    null;
    r6843 := (r6842);
    r6844 := "0";
    null;
    r6845 := (r6844);
    r6846 := "1";
    null;
    r6847 := (r6846);
    r6848 := "1";
    null;
    r6849 := (r6848);
    r6850 := "0";
    null;
    r6851 := (r6850);
    r6852 := "0";
    null;
    r6853 := (r6852);
    r6854 := "0";
    null;
    r6855 := (r6854);
    r6856 := "1";
    null;
    r6857 := (r6856);
    r6858 := "1";
    null;
    r6859 := (r6858);
    r6860 := "0";
    null;
    r6861 := (r6860);
    r6862 := "1";
    null;
    r6863 := (r6862);
    r6864 := "1";
    null;
    r6865 := (r6864);
    r6866 := "0";
    null;
    r6867 := (r6866);
    r6868 := "1";
    null;
    r6869 := (r6868);
    r6870 := "1";
    null;
    r6871 := (r6870);
    r6872 := "1";
    null;
    r6873 := (r6872);
    r6874 := "1";
    null;
    r6875 := (r6874);
    r6811 := (r6813 & r6815 & r6817 & r6819 & r6821 & r6823 & r6825 & r6827 & r6829 & r6831 & r6833 & r6835 & r6837 & r6839 & r6841 & r6843 & r6845 & r6847 & r6849 & r6851 & r6853 & r6855 & r6857 & r6859 & r6861 & r6863 & r6865 & r6867 & r6869 & r6871 & r6873 & r6875);
    return r6811;
  end rewire_MetaprogrammingRWw78a5636f_6810;
  function rewire_MetaprogrammingRWw748f82ee_6741 return std_logic_vector
  is
    variable r6806 : std_logic_vector(0 to 0) := (others => '0');
    variable r6805 : std_logic_vector(0 to 0) := (others => '0');
    variable r6804 : std_logic_vector(0 to 0) := (others => '0');
    variable r6803 : std_logic_vector(0 to 0) := (others => '0');
    variable r6802 : std_logic_vector(0 to 0) := (others => '0');
    variable r6801 : std_logic_vector(0 to 0) := (others => '0');
    variable r6800 : std_logic_vector(0 to 0) := (others => '0');
    variable r6799 : std_logic_vector(0 to 0) := (others => '0');
    variable r6798 : std_logic_vector(0 to 0) := (others => '0');
    variable r6797 : std_logic_vector(0 to 0) := (others => '0');
    variable r6796 : std_logic_vector(0 to 0) := (others => '0');
    variable r6795 : std_logic_vector(0 to 0) := (others => '0');
    variable r6794 : std_logic_vector(0 to 0) := (others => '0');
    variable r6793 : std_logic_vector(0 to 0) := (others => '0');
    variable r6792 : std_logic_vector(0 to 0) := (others => '0');
    variable r6791 : std_logic_vector(0 to 0) := (others => '0');
    variable r6790 : std_logic_vector(0 to 0) := (others => '0');
    variable r6789 : std_logic_vector(0 to 0) := (others => '0');
    variable r6788 : std_logic_vector(0 to 0) := (others => '0');
    variable r6787 : std_logic_vector(0 to 0) := (others => '0');
    variable r6786 : std_logic_vector(0 to 0) := (others => '0');
    variable r6785 : std_logic_vector(0 to 0) := (others => '0');
    variable r6784 : std_logic_vector(0 to 0) := (others => '0');
    variable r6783 : std_logic_vector(0 to 0) := (others => '0');
    variable r6782 : std_logic_vector(0 to 0) := (others => '0');
    variable r6781 : std_logic_vector(0 to 0) := (others => '0');
    variable r6780 : std_logic_vector(0 to 0) := (others => '0');
    variable r6779 : std_logic_vector(0 to 0) := (others => '0');
    variable r6778 : std_logic_vector(0 to 0) := (others => '0');
    variable r6777 : std_logic_vector(0 to 0) := (others => '0');
    variable r6776 : std_logic_vector(0 to 0) := (others => '0');
    variable r6775 : std_logic_vector(0 to 0) := (others => '0');
    variable r6774 : std_logic_vector(0 to 0) := (others => '0');
    variable r6773 : std_logic_vector(0 to 0) := (others => '0');
    variable r6772 : std_logic_vector(0 to 0) := (others => '0');
    variable r6771 : std_logic_vector(0 to 0) := (others => '0');
    variable r6770 : std_logic_vector(0 to 0) := (others => '0');
    variable r6769 : std_logic_vector(0 to 0) := (others => '0');
    variable r6768 : std_logic_vector(0 to 0) := (others => '0');
    variable r6767 : std_logic_vector(0 to 0) := (others => '0');
    variable r6766 : std_logic_vector(0 to 0) := (others => '0');
    variable r6765 : std_logic_vector(0 to 0) := (others => '0');
    variable r6764 : std_logic_vector(0 to 0) := (others => '0');
    variable r6763 : std_logic_vector(0 to 0) := (others => '0');
    variable r6762 : std_logic_vector(0 to 0) := (others => '0');
    variable r6761 : std_logic_vector(0 to 0) := (others => '0');
    variable r6760 : std_logic_vector(0 to 0) := (others => '0');
    variable r6759 : std_logic_vector(0 to 0) := (others => '0');
    variable r6758 : std_logic_vector(0 to 0) := (others => '0');
    variable r6757 : std_logic_vector(0 to 0) := (others => '0');
    variable r6756 : std_logic_vector(0 to 0) := (others => '0');
    variable r6755 : std_logic_vector(0 to 0) := (others => '0');
    variable r6754 : std_logic_vector(0 to 0) := (others => '0');
    variable r6753 : std_logic_vector(0 to 0) := (others => '0');
    variable r6752 : std_logic_vector(0 to 0) := (others => '0');
    variable r6751 : std_logic_vector(0 to 0) := (others => '0');
    variable r6750 : std_logic_vector(0 to 0) := (others => '0');
    variable r6749 : std_logic_vector(0 to 0) := (others => '0');
    variable r6748 : std_logic_vector(0 to 0) := (others => '0');
    variable r6747 : std_logic_vector(0 to 0) := (others => '0');
    variable r6746 : std_logic_vector(0 to 0) := (others => '0');
    variable r6745 : std_logic_vector(0 to 0) := (others => '0');
    variable r6744 : std_logic_vector(0 to 0) := (others => '0');
    variable r6743 : std_logic_vector(0 to 0) := (others => '0');
    variable r6742 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r6743 := "0";
    null;
    r6744 := (r6743);
    r6745 := "1";
    null;
    r6746 := (r6745);
    r6747 := "1";
    null;
    r6748 := (r6747);
    r6749 := "1";
    null;
    r6750 := (r6749);
    r6751 := "0";
    null;
    r6752 := (r6751);
    r6753 := "1";
    null;
    r6754 := (r6753);
    r6755 := "0";
    null;
    r6756 := (r6755);
    r6757 := "0";
    null;
    r6758 := (r6757);
    r6759 := "1";
    null;
    r6760 := (r6759);
    r6761 := "0";
    null;
    r6762 := (r6761);
    r6763 := "0";
    null;
    r6764 := (r6763);
    r6765 := "0";
    null;
    r6766 := (r6765);
    r6767 := "1";
    null;
    r6768 := (r6767);
    r6769 := "1";
    null;
    r6770 := (r6769);
    r6771 := "1";
    null;
    r6772 := (r6771);
    r6773 := "1";
    null;
    r6774 := (r6773);
    r6775 := "1";
    null;
    r6776 := (r6775);
    r6777 := "0";
    null;
    r6778 := (r6777);
    r6779 := "0";
    null;
    r6780 := (r6779);
    r6781 := "0";
    null;
    r6782 := (r6781);
    r6783 := "0";
    null;
    r6784 := (r6783);
    r6785 := "0";
    null;
    r6786 := (r6785);
    r6787 := "1";
    null;
    r6788 := (r6787);
    r6789 := "0";
    null;
    r6790 := (r6789);
    r6791 := "1";
    null;
    r6792 := (r6791);
    r6793 := "1";
    null;
    r6794 := (r6793);
    r6795 := "1";
    null;
    r6796 := (r6795);
    r6797 := "0";
    null;
    r6798 := (r6797);
    r6799 := "1";
    null;
    r6800 := (r6799);
    r6801 := "1";
    null;
    r6802 := (r6801);
    r6803 := "1";
    null;
    r6804 := (r6803);
    r6805 := "0";
    null;
    r6806 := (r6805);
    r6742 := (r6744 & r6746 & r6748 & r6750 & r6752 & r6754 & r6756 & r6758 & r6760 & r6762 & r6764 & r6766 & r6768 & r6770 & r6772 & r6774 & r6776 & r6778 & r6780 & r6782 & r6784 & r6786 & r6788 & r6790 & r6792 & r6794 & r6796 & r6798 & r6800 & r6802 & r6804 & r6806);
    return r6742;
  end rewire_MetaprogrammingRWw748f82ee_6741;
  function rewire_MetaprogrammingRWw682e6ff3_6672 return std_logic_vector
  is
    variable r6737 : std_logic_vector(0 to 0) := (others => '0');
    variable r6736 : std_logic_vector(0 to 0) := (others => '0');
    variable r6735 : std_logic_vector(0 to 0) := (others => '0');
    variable r6734 : std_logic_vector(0 to 0) := (others => '0');
    variable r6733 : std_logic_vector(0 to 0) := (others => '0');
    variable r6732 : std_logic_vector(0 to 0) := (others => '0');
    variable r6731 : std_logic_vector(0 to 0) := (others => '0');
    variable r6730 : std_logic_vector(0 to 0) := (others => '0');
    variable r6729 : std_logic_vector(0 to 0) := (others => '0');
    variable r6728 : std_logic_vector(0 to 0) := (others => '0');
    variable r6727 : std_logic_vector(0 to 0) := (others => '0');
    variable r6726 : std_logic_vector(0 to 0) := (others => '0');
    variable r6725 : std_logic_vector(0 to 0) := (others => '0');
    variable r6724 : std_logic_vector(0 to 0) := (others => '0');
    variable r6723 : std_logic_vector(0 to 0) := (others => '0');
    variable r6722 : std_logic_vector(0 to 0) := (others => '0');
    variable r6721 : std_logic_vector(0 to 0) := (others => '0');
    variable r6720 : std_logic_vector(0 to 0) := (others => '0');
    variable r6719 : std_logic_vector(0 to 0) := (others => '0');
    variable r6718 : std_logic_vector(0 to 0) := (others => '0');
    variable r6717 : std_logic_vector(0 to 0) := (others => '0');
    variable r6716 : std_logic_vector(0 to 0) := (others => '0');
    variable r6715 : std_logic_vector(0 to 0) := (others => '0');
    variable r6714 : std_logic_vector(0 to 0) := (others => '0');
    variable r6713 : std_logic_vector(0 to 0) := (others => '0');
    variable r6712 : std_logic_vector(0 to 0) := (others => '0');
    variable r6711 : std_logic_vector(0 to 0) := (others => '0');
    variable r6710 : std_logic_vector(0 to 0) := (others => '0');
    variable r6709 : std_logic_vector(0 to 0) := (others => '0');
    variable r6708 : std_logic_vector(0 to 0) := (others => '0');
    variable r6707 : std_logic_vector(0 to 0) := (others => '0');
    variable r6706 : std_logic_vector(0 to 0) := (others => '0');
    variable r6705 : std_logic_vector(0 to 0) := (others => '0');
    variable r6704 : std_logic_vector(0 to 0) := (others => '0');
    variable r6703 : std_logic_vector(0 to 0) := (others => '0');
    variable r6702 : std_logic_vector(0 to 0) := (others => '0');
    variable r6701 : std_logic_vector(0 to 0) := (others => '0');
    variable r6700 : std_logic_vector(0 to 0) := (others => '0');
    variable r6699 : std_logic_vector(0 to 0) := (others => '0');
    variable r6698 : std_logic_vector(0 to 0) := (others => '0');
    variable r6697 : std_logic_vector(0 to 0) := (others => '0');
    variable r6696 : std_logic_vector(0 to 0) := (others => '0');
    variable r6695 : std_logic_vector(0 to 0) := (others => '0');
    variable r6694 : std_logic_vector(0 to 0) := (others => '0');
    variable r6693 : std_logic_vector(0 to 0) := (others => '0');
    variable r6692 : std_logic_vector(0 to 0) := (others => '0');
    variable r6691 : std_logic_vector(0 to 0) := (others => '0');
    variable r6690 : std_logic_vector(0 to 0) := (others => '0');
    variable r6689 : std_logic_vector(0 to 0) := (others => '0');
    variable r6688 : std_logic_vector(0 to 0) := (others => '0');
    variable r6687 : std_logic_vector(0 to 0) := (others => '0');
    variable r6686 : std_logic_vector(0 to 0) := (others => '0');
    variable r6685 : std_logic_vector(0 to 0) := (others => '0');
    variable r6684 : std_logic_vector(0 to 0) := (others => '0');
    variable r6683 : std_logic_vector(0 to 0) := (others => '0');
    variable r6682 : std_logic_vector(0 to 0) := (others => '0');
    variable r6681 : std_logic_vector(0 to 0) := (others => '0');
    variable r6680 : std_logic_vector(0 to 0) := (others => '0');
    variable r6679 : std_logic_vector(0 to 0) := (others => '0');
    variable r6678 : std_logic_vector(0 to 0) := (others => '0');
    variable r6677 : std_logic_vector(0 to 0) := (others => '0');
    variable r6676 : std_logic_vector(0 to 0) := (others => '0');
    variable r6675 : std_logic_vector(0 to 0) := (others => '0');
    variable r6674 : std_logic_vector(0 to 0) := (others => '0');
    variable r6673 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r6674 := "0";
    null;
    r6675 := (r6674);
    r6676 := "1";
    null;
    r6677 := (r6676);
    r6678 := "1";
    null;
    r6679 := (r6678);
    r6680 := "0";
    null;
    r6681 := (r6680);
    r6682 := "1";
    null;
    r6683 := (r6682);
    r6684 := "0";
    null;
    r6685 := (r6684);
    r6686 := "0";
    null;
    r6687 := (r6686);
    r6688 := "0";
    null;
    r6689 := (r6688);
    r6690 := "0";
    null;
    r6691 := (r6690);
    r6692 := "0";
    null;
    r6693 := (r6692);
    r6694 := "1";
    null;
    r6695 := (r6694);
    r6696 := "0";
    null;
    r6697 := (r6696);
    r6698 := "1";
    null;
    r6699 := (r6698);
    r6700 := "1";
    null;
    r6701 := (r6700);
    r6702 := "1";
    null;
    r6703 := (r6702);
    r6704 := "0";
    null;
    r6705 := (r6704);
    r6706 := "0";
    null;
    r6707 := (r6706);
    r6708 := "1";
    null;
    r6709 := (r6708);
    r6710 := "1";
    null;
    r6711 := (r6710);
    r6712 := "0";
    null;
    r6713 := (r6712);
    r6714 := "1";
    null;
    r6715 := (r6714);
    r6716 := "1";
    null;
    r6717 := (r6716);
    r6718 := "1";
    null;
    r6719 := (r6718);
    r6720 := "1";
    null;
    r6721 := (r6720);
    r6722 := "1";
    null;
    r6723 := (r6722);
    r6724 := "1";
    null;
    r6725 := (r6724);
    r6726 := "1";
    null;
    r6727 := (r6726);
    r6728 := "1";
    null;
    r6729 := (r6728);
    r6730 := "0";
    null;
    r6731 := (r6730);
    r6732 := "0";
    null;
    r6733 := (r6732);
    r6734 := "1";
    null;
    r6735 := (r6734);
    r6736 := "1";
    null;
    r6737 := (r6736);
    r6673 := (r6675 & r6677 & r6679 & r6681 & r6683 & r6685 & r6687 & r6689 & r6691 & r6693 & r6695 & r6697 & r6699 & r6701 & r6703 & r6705 & r6707 & r6709 & r6711 & r6713 & r6715 & r6717 & r6719 & r6721 & r6723 & r6725 & r6727 & r6729 & r6731 & r6733 & r6735 & r6737);
    return r6673;
  end rewire_MetaprogrammingRWw682e6ff3_6672;
  function rewire_MetaprogrammingRWw5b9cca4f_6603 return std_logic_vector
  is
    variable r6668 : std_logic_vector(0 to 0) := (others => '0');
    variable r6667 : std_logic_vector(0 to 0) := (others => '0');
    variable r6666 : std_logic_vector(0 to 0) := (others => '0');
    variable r6665 : std_logic_vector(0 to 0) := (others => '0');
    variable r6664 : std_logic_vector(0 to 0) := (others => '0');
    variable r6663 : std_logic_vector(0 to 0) := (others => '0');
    variable r6662 : std_logic_vector(0 to 0) := (others => '0');
    variable r6661 : std_logic_vector(0 to 0) := (others => '0');
    variable r6660 : std_logic_vector(0 to 0) := (others => '0');
    variable r6659 : std_logic_vector(0 to 0) := (others => '0');
    variable r6658 : std_logic_vector(0 to 0) := (others => '0');
    variable r6657 : std_logic_vector(0 to 0) := (others => '0');
    variable r6656 : std_logic_vector(0 to 0) := (others => '0');
    variable r6655 : std_logic_vector(0 to 0) := (others => '0');
    variable r6654 : std_logic_vector(0 to 0) := (others => '0');
    variable r6653 : std_logic_vector(0 to 0) := (others => '0');
    variable r6652 : std_logic_vector(0 to 0) := (others => '0');
    variable r6651 : std_logic_vector(0 to 0) := (others => '0');
    variable r6650 : std_logic_vector(0 to 0) := (others => '0');
    variable r6649 : std_logic_vector(0 to 0) := (others => '0');
    variable r6648 : std_logic_vector(0 to 0) := (others => '0');
    variable r6647 : std_logic_vector(0 to 0) := (others => '0');
    variable r6646 : std_logic_vector(0 to 0) := (others => '0');
    variable r6645 : std_logic_vector(0 to 0) := (others => '0');
    variable r6644 : std_logic_vector(0 to 0) := (others => '0');
    variable r6643 : std_logic_vector(0 to 0) := (others => '0');
    variable r6642 : std_logic_vector(0 to 0) := (others => '0');
    variable r6641 : std_logic_vector(0 to 0) := (others => '0');
    variable r6640 : std_logic_vector(0 to 0) := (others => '0');
    variable r6639 : std_logic_vector(0 to 0) := (others => '0');
    variable r6638 : std_logic_vector(0 to 0) := (others => '0');
    variable r6637 : std_logic_vector(0 to 0) := (others => '0');
    variable r6636 : std_logic_vector(0 to 0) := (others => '0');
    variable r6635 : std_logic_vector(0 to 0) := (others => '0');
    variable r6634 : std_logic_vector(0 to 0) := (others => '0');
    variable r6633 : std_logic_vector(0 to 0) := (others => '0');
    variable r6632 : std_logic_vector(0 to 0) := (others => '0');
    variable r6631 : std_logic_vector(0 to 0) := (others => '0');
    variable r6630 : std_logic_vector(0 to 0) := (others => '0');
    variable r6629 : std_logic_vector(0 to 0) := (others => '0');
    variable r6628 : std_logic_vector(0 to 0) := (others => '0');
    variable r6627 : std_logic_vector(0 to 0) := (others => '0');
    variable r6626 : std_logic_vector(0 to 0) := (others => '0');
    variable r6625 : std_logic_vector(0 to 0) := (others => '0');
    variable r6624 : std_logic_vector(0 to 0) := (others => '0');
    variable r6623 : std_logic_vector(0 to 0) := (others => '0');
    variable r6622 : std_logic_vector(0 to 0) := (others => '0');
    variable r6621 : std_logic_vector(0 to 0) := (others => '0');
    variable r6620 : std_logic_vector(0 to 0) := (others => '0');
    variable r6619 : std_logic_vector(0 to 0) := (others => '0');
    variable r6618 : std_logic_vector(0 to 0) := (others => '0');
    variable r6617 : std_logic_vector(0 to 0) := (others => '0');
    variable r6616 : std_logic_vector(0 to 0) := (others => '0');
    variable r6615 : std_logic_vector(0 to 0) := (others => '0');
    variable r6614 : std_logic_vector(0 to 0) := (others => '0');
    variable r6613 : std_logic_vector(0 to 0) := (others => '0');
    variable r6612 : std_logic_vector(0 to 0) := (others => '0');
    variable r6611 : std_logic_vector(0 to 0) := (others => '0');
    variable r6610 : std_logic_vector(0 to 0) := (others => '0');
    variable r6609 : std_logic_vector(0 to 0) := (others => '0');
    variable r6608 : std_logic_vector(0 to 0) := (others => '0');
    variable r6607 : std_logic_vector(0 to 0) := (others => '0');
    variable r6606 : std_logic_vector(0 to 0) := (others => '0');
    variable r6605 : std_logic_vector(0 to 0) := (others => '0');
    variable r6604 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r6605 := "0";
    null;
    r6606 := (r6605);
    r6607 := "1";
    null;
    r6608 := (r6607);
    r6609 := "0";
    null;
    r6610 := (r6609);
    r6611 := "1";
    null;
    r6612 := (r6611);
    r6613 := "1";
    null;
    r6614 := (r6613);
    r6615 := "0";
    null;
    r6616 := (r6615);
    r6617 := "1";
    null;
    r6618 := (r6617);
    r6619 := "1";
    null;
    r6620 := (r6619);
    r6621 := "1";
    null;
    r6622 := (r6621);
    r6623 := "0";
    null;
    r6624 := (r6623);
    r6625 := "0";
    null;
    r6626 := (r6625);
    r6627 := "1";
    null;
    r6628 := (r6627);
    r6629 := "1";
    null;
    r6630 := (r6629);
    r6631 := "1";
    null;
    r6632 := (r6631);
    r6633 := "0";
    null;
    r6634 := (r6633);
    r6635 := "0";
    null;
    r6636 := (r6635);
    r6637 := "1";
    null;
    r6638 := (r6637);
    r6639 := "1";
    null;
    r6640 := (r6639);
    r6641 := "0";
    null;
    r6642 := (r6641);
    r6643 := "0";
    null;
    r6644 := (r6643);
    r6645 := "1";
    null;
    r6646 := (r6645);
    r6647 := "0";
    null;
    r6648 := (r6647);
    r6649 := "1";
    null;
    r6650 := (r6649);
    r6651 := "0";
    null;
    r6652 := (r6651);
    r6653 := "0";
    null;
    r6654 := (r6653);
    r6655 := "1";
    null;
    r6656 := (r6655);
    r6657 := "0";
    null;
    r6658 := (r6657);
    r6659 := "0";
    null;
    r6660 := (r6659);
    r6661 := "1";
    null;
    r6662 := (r6661);
    r6663 := "1";
    null;
    r6664 := (r6663);
    r6665 := "1";
    null;
    r6666 := (r6665);
    r6667 := "1";
    null;
    r6668 := (r6667);
    r6604 := (r6606 & r6608 & r6610 & r6612 & r6614 & r6616 & r6618 & r6620 & r6622 & r6624 & r6626 & r6628 & r6630 & r6632 & r6634 & r6636 & r6638 & r6640 & r6642 & r6644 & r6646 & r6648 & r6650 & r6652 & r6654 & r6656 & r6658 & r6660 & r6662 & r6664 & r6666 & r6668);
    return r6604;
  end rewire_MetaprogrammingRWw5b9cca4f_6603;
  function rewire_MetaprogrammingRWw4ed8aa4a_6534 return std_logic_vector
  is
    variable r6599 : std_logic_vector(0 to 0) := (others => '0');
    variable r6598 : std_logic_vector(0 to 0) := (others => '0');
    variable r6597 : std_logic_vector(0 to 0) := (others => '0');
    variable r6596 : std_logic_vector(0 to 0) := (others => '0');
    variable r6595 : std_logic_vector(0 to 0) := (others => '0');
    variable r6594 : std_logic_vector(0 to 0) := (others => '0');
    variable r6593 : std_logic_vector(0 to 0) := (others => '0');
    variable r6592 : std_logic_vector(0 to 0) := (others => '0');
    variable r6591 : std_logic_vector(0 to 0) := (others => '0');
    variable r6590 : std_logic_vector(0 to 0) := (others => '0');
    variable r6589 : std_logic_vector(0 to 0) := (others => '0');
    variable r6588 : std_logic_vector(0 to 0) := (others => '0');
    variable r6587 : std_logic_vector(0 to 0) := (others => '0');
    variable r6586 : std_logic_vector(0 to 0) := (others => '0');
    variable r6585 : std_logic_vector(0 to 0) := (others => '0');
    variable r6584 : std_logic_vector(0 to 0) := (others => '0');
    variable r6583 : std_logic_vector(0 to 0) := (others => '0');
    variable r6582 : std_logic_vector(0 to 0) := (others => '0');
    variable r6581 : std_logic_vector(0 to 0) := (others => '0');
    variable r6580 : std_logic_vector(0 to 0) := (others => '0');
    variable r6579 : std_logic_vector(0 to 0) := (others => '0');
    variable r6578 : std_logic_vector(0 to 0) := (others => '0');
    variable r6577 : std_logic_vector(0 to 0) := (others => '0');
    variable r6576 : std_logic_vector(0 to 0) := (others => '0');
    variable r6575 : std_logic_vector(0 to 0) := (others => '0');
    variable r6574 : std_logic_vector(0 to 0) := (others => '0');
    variable r6573 : std_logic_vector(0 to 0) := (others => '0');
    variable r6572 : std_logic_vector(0 to 0) := (others => '0');
    variable r6571 : std_logic_vector(0 to 0) := (others => '0');
    variable r6570 : std_logic_vector(0 to 0) := (others => '0');
    variable r6569 : std_logic_vector(0 to 0) := (others => '0');
    variable r6568 : std_logic_vector(0 to 0) := (others => '0');
    variable r6567 : std_logic_vector(0 to 0) := (others => '0');
    variable r6566 : std_logic_vector(0 to 0) := (others => '0');
    variable r6565 : std_logic_vector(0 to 0) := (others => '0');
    variable r6564 : std_logic_vector(0 to 0) := (others => '0');
    variable r6563 : std_logic_vector(0 to 0) := (others => '0');
    variable r6562 : std_logic_vector(0 to 0) := (others => '0');
    variable r6561 : std_logic_vector(0 to 0) := (others => '0');
    variable r6560 : std_logic_vector(0 to 0) := (others => '0');
    variable r6559 : std_logic_vector(0 to 0) := (others => '0');
    variable r6558 : std_logic_vector(0 to 0) := (others => '0');
    variable r6557 : std_logic_vector(0 to 0) := (others => '0');
    variable r6556 : std_logic_vector(0 to 0) := (others => '0');
    variable r6555 : std_logic_vector(0 to 0) := (others => '0');
    variable r6554 : std_logic_vector(0 to 0) := (others => '0');
    variable r6553 : std_logic_vector(0 to 0) := (others => '0');
    variable r6552 : std_logic_vector(0 to 0) := (others => '0');
    variable r6551 : std_logic_vector(0 to 0) := (others => '0');
    variable r6550 : std_logic_vector(0 to 0) := (others => '0');
    variable r6549 : std_logic_vector(0 to 0) := (others => '0');
    variable r6548 : std_logic_vector(0 to 0) := (others => '0');
    variable r6547 : std_logic_vector(0 to 0) := (others => '0');
    variable r6546 : std_logic_vector(0 to 0) := (others => '0');
    variable r6545 : std_logic_vector(0 to 0) := (others => '0');
    variable r6544 : std_logic_vector(0 to 0) := (others => '0');
    variable r6543 : std_logic_vector(0 to 0) := (others => '0');
    variable r6542 : std_logic_vector(0 to 0) := (others => '0');
    variable r6541 : std_logic_vector(0 to 0) := (others => '0');
    variable r6540 : std_logic_vector(0 to 0) := (others => '0');
    variable r6539 : std_logic_vector(0 to 0) := (others => '0');
    variable r6538 : std_logic_vector(0 to 0) := (others => '0');
    variable r6537 : std_logic_vector(0 to 0) := (others => '0');
    variable r6536 : std_logic_vector(0 to 0) := (others => '0');
    variable r6535 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r6536 := "0";
    null;
    r6537 := (r6536);
    r6538 := "1";
    null;
    r6539 := (r6538);
    r6540 := "0";
    null;
    r6541 := (r6540);
    r6542 := "0";
    null;
    r6543 := (r6542);
    r6544 := "1";
    null;
    r6545 := (r6544);
    r6546 := "1";
    null;
    r6547 := (r6546);
    r6548 := "1";
    null;
    r6549 := (r6548);
    r6550 := "0";
    null;
    r6551 := (r6550);
    r6552 := "1";
    null;
    r6553 := (r6552);
    r6554 := "1";
    null;
    r6555 := (r6554);
    r6556 := "0";
    null;
    r6557 := (r6556);
    r6558 := "1";
    null;
    r6559 := (r6558);
    r6560 := "1";
    null;
    r6561 := (r6560);
    r6562 := "0";
    null;
    r6563 := (r6562);
    r6564 := "0";
    null;
    r6565 := (r6564);
    r6566 := "0";
    null;
    r6567 := (r6566);
    r6568 := "1";
    null;
    r6569 := (r6568);
    r6570 := "0";
    null;
    r6571 := (r6570);
    r6572 := "1";
    null;
    r6573 := (r6572);
    r6574 := "0";
    null;
    r6575 := (r6574);
    r6576 := "1";
    null;
    r6577 := (r6576);
    r6578 := "0";
    null;
    r6579 := (r6578);
    r6580 := "1";
    null;
    r6581 := (r6580);
    r6582 := "0";
    null;
    r6583 := (r6582);
    r6584 := "0";
    null;
    r6585 := (r6584);
    r6586 := "1";
    null;
    r6587 := (r6586);
    r6588 := "0";
    null;
    r6589 := (r6588);
    r6590 := "0";
    null;
    r6591 := (r6590);
    r6592 := "1";
    null;
    r6593 := (r6592);
    r6594 := "0";
    null;
    r6595 := (r6594);
    r6596 := "1";
    null;
    r6597 := (r6596);
    r6598 := "0";
    null;
    r6599 := (r6598);
    r6535 := (r6537 & r6539 & r6541 & r6543 & r6545 & r6547 & r6549 & r6551 & r6553 & r6555 & r6557 & r6559 & r6561 & r6563 & r6565 & r6567 & r6569 & r6571 & r6573 & r6575 & r6577 & r6579 & r6581 & r6583 & r6585 & r6587 & r6589 & r6591 & r6593 & r6595 & r6597 & r6599);
    return r6535;
  end rewire_MetaprogrammingRWw4ed8aa4a_6534;
  function rewire_MetaprogrammingRWw391c0cb3_6465 return std_logic_vector
  is
    variable r6530 : std_logic_vector(0 to 0) := (others => '0');
    variable r6529 : std_logic_vector(0 to 0) := (others => '0');
    variable r6528 : std_logic_vector(0 to 0) := (others => '0');
    variable r6527 : std_logic_vector(0 to 0) := (others => '0');
    variable r6526 : std_logic_vector(0 to 0) := (others => '0');
    variable r6525 : std_logic_vector(0 to 0) := (others => '0');
    variable r6524 : std_logic_vector(0 to 0) := (others => '0');
    variable r6523 : std_logic_vector(0 to 0) := (others => '0');
    variable r6522 : std_logic_vector(0 to 0) := (others => '0');
    variable r6521 : std_logic_vector(0 to 0) := (others => '0');
    variable r6520 : std_logic_vector(0 to 0) := (others => '0');
    variable r6519 : std_logic_vector(0 to 0) := (others => '0');
    variable r6518 : std_logic_vector(0 to 0) := (others => '0');
    variable r6517 : std_logic_vector(0 to 0) := (others => '0');
    variable r6516 : std_logic_vector(0 to 0) := (others => '0');
    variable r6515 : std_logic_vector(0 to 0) := (others => '0');
    variable r6514 : std_logic_vector(0 to 0) := (others => '0');
    variable r6513 : std_logic_vector(0 to 0) := (others => '0');
    variable r6512 : std_logic_vector(0 to 0) := (others => '0');
    variable r6511 : std_logic_vector(0 to 0) := (others => '0');
    variable r6510 : std_logic_vector(0 to 0) := (others => '0');
    variable r6509 : std_logic_vector(0 to 0) := (others => '0');
    variable r6508 : std_logic_vector(0 to 0) := (others => '0');
    variable r6507 : std_logic_vector(0 to 0) := (others => '0');
    variable r6506 : std_logic_vector(0 to 0) := (others => '0');
    variable r6505 : std_logic_vector(0 to 0) := (others => '0');
    variable r6504 : std_logic_vector(0 to 0) := (others => '0');
    variable r6503 : std_logic_vector(0 to 0) := (others => '0');
    variable r6502 : std_logic_vector(0 to 0) := (others => '0');
    variable r6501 : std_logic_vector(0 to 0) := (others => '0');
    variable r6500 : std_logic_vector(0 to 0) := (others => '0');
    variable r6499 : std_logic_vector(0 to 0) := (others => '0');
    variable r6498 : std_logic_vector(0 to 0) := (others => '0');
    variable r6497 : std_logic_vector(0 to 0) := (others => '0');
    variable r6496 : std_logic_vector(0 to 0) := (others => '0');
    variable r6495 : std_logic_vector(0 to 0) := (others => '0');
    variable r6494 : std_logic_vector(0 to 0) := (others => '0');
    variable r6493 : std_logic_vector(0 to 0) := (others => '0');
    variable r6492 : std_logic_vector(0 to 0) := (others => '0');
    variable r6491 : std_logic_vector(0 to 0) := (others => '0');
    variable r6490 : std_logic_vector(0 to 0) := (others => '0');
    variable r6489 : std_logic_vector(0 to 0) := (others => '0');
    variable r6488 : std_logic_vector(0 to 0) := (others => '0');
    variable r6487 : std_logic_vector(0 to 0) := (others => '0');
    variable r6486 : std_logic_vector(0 to 0) := (others => '0');
    variable r6485 : std_logic_vector(0 to 0) := (others => '0');
    variable r6484 : std_logic_vector(0 to 0) := (others => '0');
    variable r6483 : std_logic_vector(0 to 0) := (others => '0');
    variable r6482 : std_logic_vector(0 to 0) := (others => '0');
    variable r6481 : std_logic_vector(0 to 0) := (others => '0');
    variable r6480 : std_logic_vector(0 to 0) := (others => '0');
    variable r6479 : std_logic_vector(0 to 0) := (others => '0');
    variable r6478 : std_logic_vector(0 to 0) := (others => '0');
    variable r6477 : std_logic_vector(0 to 0) := (others => '0');
    variable r6476 : std_logic_vector(0 to 0) := (others => '0');
    variable r6475 : std_logic_vector(0 to 0) := (others => '0');
    variable r6474 : std_logic_vector(0 to 0) := (others => '0');
    variable r6473 : std_logic_vector(0 to 0) := (others => '0');
    variable r6472 : std_logic_vector(0 to 0) := (others => '0');
    variable r6471 : std_logic_vector(0 to 0) := (others => '0');
    variable r6470 : std_logic_vector(0 to 0) := (others => '0');
    variable r6469 : std_logic_vector(0 to 0) := (others => '0');
    variable r6468 : std_logic_vector(0 to 0) := (others => '0');
    variable r6467 : std_logic_vector(0 to 0) := (others => '0');
    variable r6466 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r6467 := "0";
    null;
    r6468 := (r6467);
    r6469 := "0";
    null;
    r6470 := (r6469);
    r6471 := "1";
    null;
    r6472 := (r6471);
    r6473 := "1";
    null;
    r6474 := (r6473);
    r6475 := "1";
    null;
    r6476 := (r6475);
    r6477 := "0";
    null;
    r6478 := (r6477);
    r6479 := "0";
    null;
    r6480 := (r6479);
    r6481 := "1";
    null;
    r6482 := (r6481);
    r6483 := "0";
    null;
    r6484 := (r6483);
    r6485 := "0";
    null;
    r6486 := (r6485);
    r6487 := "0";
    null;
    r6488 := (r6487);
    r6489 := "1";
    null;
    r6490 := (r6489);
    r6491 := "1";
    null;
    r6492 := (r6491);
    r6493 := "1";
    null;
    r6494 := (r6493);
    r6495 := "0";
    null;
    r6496 := (r6495);
    r6497 := "0";
    null;
    r6498 := (r6497);
    r6499 := "0";
    null;
    r6500 := (r6499);
    r6501 := "0";
    null;
    r6502 := (r6501);
    r6503 := "0";
    null;
    r6504 := (r6503);
    r6505 := "0";
    null;
    r6506 := (r6505);
    r6507 := "1";
    null;
    r6508 := (r6507);
    r6509 := "1";
    null;
    r6510 := (r6509);
    r6511 := "0";
    null;
    r6512 := (r6511);
    r6513 := "0";
    null;
    r6514 := (r6513);
    r6515 := "1";
    null;
    r6516 := (r6515);
    r6517 := "0";
    null;
    r6518 := (r6517);
    r6519 := "1";
    null;
    r6520 := (r6519);
    r6521 := "1";
    null;
    r6522 := (r6521);
    r6523 := "0";
    null;
    r6524 := (r6523);
    r6525 := "0";
    null;
    r6526 := (r6525);
    r6527 := "1";
    null;
    r6528 := (r6527);
    r6529 := "1";
    null;
    r6530 := (r6529);
    r6466 := (r6468 & r6470 & r6472 & r6474 & r6476 & r6478 & r6480 & r6482 & r6484 & r6486 & r6488 & r6490 & r6492 & r6494 & r6496 & r6498 & r6500 & r6502 & r6504 & r6506 & r6508 & r6510 & r6512 & r6514 & r6516 & r6518 & r6520 & r6522 & r6524 & r6526 & r6528 & r6530);
    return r6466;
  end rewire_MetaprogrammingRWw391c0cb3_6465;
  function rewire_MetaprogrammingRWw34b0bcb5_6396 return std_logic_vector
  is
    variable r6461 : std_logic_vector(0 to 0) := (others => '0');
    variable r6460 : std_logic_vector(0 to 0) := (others => '0');
    variable r6459 : std_logic_vector(0 to 0) := (others => '0');
    variable r6458 : std_logic_vector(0 to 0) := (others => '0');
    variable r6457 : std_logic_vector(0 to 0) := (others => '0');
    variable r6456 : std_logic_vector(0 to 0) := (others => '0');
    variable r6455 : std_logic_vector(0 to 0) := (others => '0');
    variable r6454 : std_logic_vector(0 to 0) := (others => '0');
    variable r6453 : std_logic_vector(0 to 0) := (others => '0');
    variable r6452 : std_logic_vector(0 to 0) := (others => '0');
    variable r6451 : std_logic_vector(0 to 0) := (others => '0');
    variable r6450 : std_logic_vector(0 to 0) := (others => '0');
    variable r6449 : std_logic_vector(0 to 0) := (others => '0');
    variable r6448 : std_logic_vector(0 to 0) := (others => '0');
    variable r6447 : std_logic_vector(0 to 0) := (others => '0');
    variable r6446 : std_logic_vector(0 to 0) := (others => '0');
    variable r6445 : std_logic_vector(0 to 0) := (others => '0');
    variable r6444 : std_logic_vector(0 to 0) := (others => '0');
    variable r6443 : std_logic_vector(0 to 0) := (others => '0');
    variable r6442 : std_logic_vector(0 to 0) := (others => '0');
    variable r6441 : std_logic_vector(0 to 0) := (others => '0');
    variable r6440 : std_logic_vector(0 to 0) := (others => '0');
    variable r6439 : std_logic_vector(0 to 0) := (others => '0');
    variable r6438 : std_logic_vector(0 to 0) := (others => '0');
    variable r6437 : std_logic_vector(0 to 0) := (others => '0');
    variable r6436 : std_logic_vector(0 to 0) := (others => '0');
    variable r6435 : std_logic_vector(0 to 0) := (others => '0');
    variable r6434 : std_logic_vector(0 to 0) := (others => '0');
    variable r6433 : std_logic_vector(0 to 0) := (others => '0');
    variable r6432 : std_logic_vector(0 to 0) := (others => '0');
    variable r6431 : std_logic_vector(0 to 0) := (others => '0');
    variable r6430 : std_logic_vector(0 to 0) := (others => '0');
    variable r6429 : std_logic_vector(0 to 0) := (others => '0');
    variable r6428 : std_logic_vector(0 to 0) := (others => '0');
    variable r6427 : std_logic_vector(0 to 0) := (others => '0');
    variable r6426 : std_logic_vector(0 to 0) := (others => '0');
    variable r6425 : std_logic_vector(0 to 0) := (others => '0');
    variable r6424 : std_logic_vector(0 to 0) := (others => '0');
    variable r6423 : std_logic_vector(0 to 0) := (others => '0');
    variable r6422 : std_logic_vector(0 to 0) := (others => '0');
    variable r6421 : std_logic_vector(0 to 0) := (others => '0');
    variable r6420 : std_logic_vector(0 to 0) := (others => '0');
    variable r6419 : std_logic_vector(0 to 0) := (others => '0');
    variable r6418 : std_logic_vector(0 to 0) := (others => '0');
    variable r6417 : std_logic_vector(0 to 0) := (others => '0');
    variable r6416 : std_logic_vector(0 to 0) := (others => '0');
    variable r6415 : std_logic_vector(0 to 0) := (others => '0');
    variable r6414 : std_logic_vector(0 to 0) := (others => '0');
    variable r6413 : std_logic_vector(0 to 0) := (others => '0');
    variable r6412 : std_logic_vector(0 to 0) := (others => '0');
    variable r6411 : std_logic_vector(0 to 0) := (others => '0');
    variable r6410 : std_logic_vector(0 to 0) := (others => '0');
    variable r6409 : std_logic_vector(0 to 0) := (others => '0');
    variable r6408 : std_logic_vector(0 to 0) := (others => '0');
    variable r6407 : std_logic_vector(0 to 0) := (others => '0');
    variable r6406 : std_logic_vector(0 to 0) := (others => '0');
    variable r6405 : std_logic_vector(0 to 0) := (others => '0');
    variable r6404 : std_logic_vector(0 to 0) := (others => '0');
    variable r6403 : std_logic_vector(0 to 0) := (others => '0');
    variable r6402 : std_logic_vector(0 to 0) := (others => '0');
    variable r6401 : std_logic_vector(0 to 0) := (others => '0');
    variable r6400 : std_logic_vector(0 to 0) := (others => '0');
    variable r6399 : std_logic_vector(0 to 0) := (others => '0');
    variable r6398 : std_logic_vector(0 to 0) := (others => '0');
    variable r6397 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r6398 := "0";
    null;
    r6399 := (r6398);
    r6400 := "0";
    null;
    r6401 := (r6400);
    r6402 := "1";
    null;
    r6403 := (r6402);
    r6404 := "1";
    null;
    r6405 := (r6404);
    r6406 := "0";
    null;
    r6407 := (r6406);
    r6408 := "1";
    null;
    r6409 := (r6408);
    r6410 := "0";
    null;
    r6411 := (r6410);
    r6412 := "0";
    null;
    r6413 := (r6412);
    r6414 := "1";
    null;
    r6415 := (r6414);
    r6416 := "0";
    null;
    r6417 := (r6416);
    r6418 := "1";
    null;
    r6419 := (r6418);
    r6420 := "1";
    null;
    r6421 := (r6420);
    r6422 := "0";
    null;
    r6423 := (r6422);
    r6424 := "0";
    null;
    r6425 := (r6424);
    r6426 := "0";
    null;
    r6427 := (r6426);
    r6428 := "0";
    null;
    r6429 := (r6428);
    r6430 := "1";
    null;
    r6431 := (r6430);
    r6432 := "0";
    null;
    r6433 := (r6432);
    r6434 := "1";
    null;
    r6435 := (r6434);
    r6436 := "1";
    null;
    r6437 := (r6436);
    r6438 := "1";
    null;
    r6439 := (r6438);
    r6440 := "1";
    null;
    r6441 := (r6440);
    r6442 := "0";
    null;
    r6443 := (r6442);
    r6444 := "0";
    null;
    r6445 := (r6444);
    r6446 := "1";
    null;
    r6447 := (r6446);
    r6448 := "0";
    null;
    r6449 := (r6448);
    r6450 := "1";
    null;
    r6451 := (r6450);
    r6452 := "1";
    null;
    r6453 := (r6452);
    r6454 := "0";
    null;
    r6455 := (r6454);
    r6456 := "1";
    null;
    r6457 := (r6456);
    r6458 := "0";
    null;
    r6459 := (r6458);
    r6460 := "1";
    null;
    r6461 := (r6460);
    r6397 := (r6399 & r6401 & r6403 & r6405 & r6407 & r6409 & r6411 & r6413 & r6415 & r6417 & r6419 & r6421 & r6423 & r6425 & r6427 & r6429 & r6431 & r6433 & r6435 & r6437 & r6439 & r6441 & r6443 & r6445 & r6447 & r6449 & r6451 & r6453 & r6455 & r6457 & r6459 & r6461);
    return r6397;
  end rewire_MetaprogrammingRWw34b0bcb5_6396;
  function rewire_MetaprogrammingRWw2748774c_6327 return std_logic_vector
  is
    variable r6392 : std_logic_vector(0 to 0) := (others => '0');
    variable r6391 : std_logic_vector(0 to 0) := (others => '0');
    variable r6390 : std_logic_vector(0 to 0) := (others => '0');
    variable r6389 : std_logic_vector(0 to 0) := (others => '0');
    variable r6388 : std_logic_vector(0 to 0) := (others => '0');
    variable r6387 : std_logic_vector(0 to 0) := (others => '0');
    variable r6386 : std_logic_vector(0 to 0) := (others => '0');
    variable r6385 : std_logic_vector(0 to 0) := (others => '0');
    variable r6384 : std_logic_vector(0 to 0) := (others => '0');
    variable r6383 : std_logic_vector(0 to 0) := (others => '0');
    variable r6382 : std_logic_vector(0 to 0) := (others => '0');
    variable r6381 : std_logic_vector(0 to 0) := (others => '0');
    variable r6380 : std_logic_vector(0 to 0) := (others => '0');
    variable r6379 : std_logic_vector(0 to 0) := (others => '0');
    variable r6378 : std_logic_vector(0 to 0) := (others => '0');
    variable r6377 : std_logic_vector(0 to 0) := (others => '0');
    variable r6376 : std_logic_vector(0 to 0) := (others => '0');
    variable r6375 : std_logic_vector(0 to 0) := (others => '0');
    variable r6374 : std_logic_vector(0 to 0) := (others => '0');
    variable r6373 : std_logic_vector(0 to 0) := (others => '0');
    variable r6372 : std_logic_vector(0 to 0) := (others => '0');
    variable r6371 : std_logic_vector(0 to 0) := (others => '0');
    variable r6370 : std_logic_vector(0 to 0) := (others => '0');
    variable r6369 : std_logic_vector(0 to 0) := (others => '0');
    variable r6368 : std_logic_vector(0 to 0) := (others => '0');
    variable r6367 : std_logic_vector(0 to 0) := (others => '0');
    variable r6366 : std_logic_vector(0 to 0) := (others => '0');
    variable r6365 : std_logic_vector(0 to 0) := (others => '0');
    variable r6364 : std_logic_vector(0 to 0) := (others => '0');
    variable r6363 : std_logic_vector(0 to 0) := (others => '0');
    variable r6362 : std_logic_vector(0 to 0) := (others => '0');
    variable r6361 : std_logic_vector(0 to 0) := (others => '0');
    variable r6360 : std_logic_vector(0 to 0) := (others => '0');
    variable r6359 : std_logic_vector(0 to 0) := (others => '0');
    variable r6358 : std_logic_vector(0 to 0) := (others => '0');
    variable r6357 : std_logic_vector(0 to 0) := (others => '0');
    variable r6356 : std_logic_vector(0 to 0) := (others => '0');
    variable r6355 : std_logic_vector(0 to 0) := (others => '0');
    variable r6354 : std_logic_vector(0 to 0) := (others => '0');
    variable r6353 : std_logic_vector(0 to 0) := (others => '0');
    variable r6352 : std_logic_vector(0 to 0) := (others => '0');
    variable r6351 : std_logic_vector(0 to 0) := (others => '0');
    variable r6350 : std_logic_vector(0 to 0) := (others => '0');
    variable r6349 : std_logic_vector(0 to 0) := (others => '0');
    variable r6348 : std_logic_vector(0 to 0) := (others => '0');
    variable r6347 : std_logic_vector(0 to 0) := (others => '0');
    variable r6346 : std_logic_vector(0 to 0) := (others => '0');
    variable r6345 : std_logic_vector(0 to 0) := (others => '0');
    variable r6344 : std_logic_vector(0 to 0) := (others => '0');
    variable r6343 : std_logic_vector(0 to 0) := (others => '0');
    variable r6342 : std_logic_vector(0 to 0) := (others => '0');
    variable r6341 : std_logic_vector(0 to 0) := (others => '0');
    variable r6340 : std_logic_vector(0 to 0) := (others => '0');
    variable r6339 : std_logic_vector(0 to 0) := (others => '0');
    variable r6338 : std_logic_vector(0 to 0) := (others => '0');
    variable r6337 : std_logic_vector(0 to 0) := (others => '0');
    variable r6336 : std_logic_vector(0 to 0) := (others => '0');
    variable r6335 : std_logic_vector(0 to 0) := (others => '0');
    variable r6334 : std_logic_vector(0 to 0) := (others => '0');
    variable r6333 : std_logic_vector(0 to 0) := (others => '0');
    variable r6332 : std_logic_vector(0 to 0) := (others => '0');
    variable r6331 : std_logic_vector(0 to 0) := (others => '0');
    variable r6330 : std_logic_vector(0 to 0) := (others => '0');
    variable r6329 : std_logic_vector(0 to 0) := (others => '0');
    variable r6328 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r6329 := "0";
    null;
    r6330 := (r6329);
    r6331 := "0";
    null;
    r6332 := (r6331);
    r6333 := "1";
    null;
    r6334 := (r6333);
    r6335 := "0";
    null;
    r6336 := (r6335);
    r6337 := "0";
    null;
    r6338 := (r6337);
    r6339 := "1";
    null;
    r6340 := (r6339);
    r6341 := "1";
    null;
    r6342 := (r6341);
    r6343 := "1";
    null;
    r6344 := (r6343);
    r6345 := "0";
    null;
    r6346 := (r6345);
    r6347 := "1";
    null;
    r6348 := (r6347);
    r6349 := "0";
    null;
    r6350 := (r6349);
    r6351 := "0";
    null;
    r6352 := (r6351);
    r6353 := "1";
    null;
    r6354 := (r6353);
    r6355 := "0";
    null;
    r6356 := (r6355);
    r6357 := "0";
    null;
    r6358 := (r6357);
    r6359 := "0";
    null;
    r6360 := (r6359);
    r6361 := "0";
    null;
    r6362 := (r6361);
    r6363 := "1";
    null;
    r6364 := (r6363);
    r6365 := "1";
    null;
    r6366 := (r6365);
    r6367 := "1";
    null;
    r6368 := (r6367);
    r6369 := "0";
    null;
    r6370 := (r6369);
    r6371 := "1";
    null;
    r6372 := (r6371);
    r6373 := "1";
    null;
    r6374 := (r6373);
    r6375 := "1";
    null;
    r6376 := (r6375);
    r6377 := "0";
    null;
    r6378 := (r6377);
    r6379 := "1";
    null;
    r6380 := (r6379);
    r6381 := "0";
    null;
    r6382 := (r6381);
    r6383 := "0";
    null;
    r6384 := (r6383);
    r6385 := "1";
    null;
    r6386 := (r6385);
    r6387 := "1";
    null;
    r6388 := (r6387);
    r6389 := "0";
    null;
    r6390 := (r6389);
    r6391 := "0";
    null;
    r6392 := (r6391);
    r6328 := (r6330 & r6332 & r6334 & r6336 & r6338 & r6340 & r6342 & r6344 & r6346 & r6348 & r6350 & r6352 & r6354 & r6356 & r6358 & r6360 & r6362 & r6364 & r6366 & r6368 & r6370 & r6372 & r6374 & r6376 & r6378 & r6380 & r6382 & r6384 & r6386 & r6388 & r6390 & r6392);
    return r6328;
  end rewire_MetaprogrammingRWw2748774c_6327;
  function rewire_MetaprogrammingRWw1e376c08_6258 return std_logic_vector
  is
    variable r6323 : std_logic_vector(0 to 0) := (others => '0');
    variable r6322 : std_logic_vector(0 to 0) := (others => '0');
    variable r6321 : std_logic_vector(0 to 0) := (others => '0');
    variable r6320 : std_logic_vector(0 to 0) := (others => '0');
    variable r6319 : std_logic_vector(0 to 0) := (others => '0');
    variable r6318 : std_logic_vector(0 to 0) := (others => '0');
    variable r6317 : std_logic_vector(0 to 0) := (others => '0');
    variable r6316 : std_logic_vector(0 to 0) := (others => '0');
    variable r6315 : std_logic_vector(0 to 0) := (others => '0');
    variable r6314 : std_logic_vector(0 to 0) := (others => '0');
    variable r6313 : std_logic_vector(0 to 0) := (others => '0');
    variable r6312 : std_logic_vector(0 to 0) := (others => '0');
    variable r6311 : std_logic_vector(0 to 0) := (others => '0');
    variable r6310 : std_logic_vector(0 to 0) := (others => '0');
    variable r6309 : std_logic_vector(0 to 0) := (others => '0');
    variable r6308 : std_logic_vector(0 to 0) := (others => '0');
    variable r6307 : std_logic_vector(0 to 0) := (others => '0');
    variable r6306 : std_logic_vector(0 to 0) := (others => '0');
    variable r6305 : std_logic_vector(0 to 0) := (others => '0');
    variable r6304 : std_logic_vector(0 to 0) := (others => '0');
    variable r6303 : std_logic_vector(0 to 0) := (others => '0');
    variable r6302 : std_logic_vector(0 to 0) := (others => '0');
    variable r6301 : std_logic_vector(0 to 0) := (others => '0');
    variable r6300 : std_logic_vector(0 to 0) := (others => '0');
    variable r6299 : std_logic_vector(0 to 0) := (others => '0');
    variable r6298 : std_logic_vector(0 to 0) := (others => '0');
    variable r6297 : std_logic_vector(0 to 0) := (others => '0');
    variable r6296 : std_logic_vector(0 to 0) := (others => '0');
    variable r6295 : std_logic_vector(0 to 0) := (others => '0');
    variable r6294 : std_logic_vector(0 to 0) := (others => '0');
    variable r6293 : std_logic_vector(0 to 0) := (others => '0');
    variable r6292 : std_logic_vector(0 to 0) := (others => '0');
    variable r6291 : std_logic_vector(0 to 0) := (others => '0');
    variable r6290 : std_logic_vector(0 to 0) := (others => '0');
    variable r6289 : std_logic_vector(0 to 0) := (others => '0');
    variable r6288 : std_logic_vector(0 to 0) := (others => '0');
    variable r6287 : std_logic_vector(0 to 0) := (others => '0');
    variable r6286 : std_logic_vector(0 to 0) := (others => '0');
    variable r6285 : std_logic_vector(0 to 0) := (others => '0');
    variable r6284 : std_logic_vector(0 to 0) := (others => '0');
    variable r6283 : std_logic_vector(0 to 0) := (others => '0');
    variable r6282 : std_logic_vector(0 to 0) := (others => '0');
    variable r6281 : std_logic_vector(0 to 0) := (others => '0');
    variable r6280 : std_logic_vector(0 to 0) := (others => '0');
    variable r6279 : std_logic_vector(0 to 0) := (others => '0');
    variable r6278 : std_logic_vector(0 to 0) := (others => '0');
    variable r6277 : std_logic_vector(0 to 0) := (others => '0');
    variable r6276 : std_logic_vector(0 to 0) := (others => '0');
    variable r6275 : std_logic_vector(0 to 0) := (others => '0');
    variable r6274 : std_logic_vector(0 to 0) := (others => '0');
    variable r6273 : std_logic_vector(0 to 0) := (others => '0');
    variable r6272 : std_logic_vector(0 to 0) := (others => '0');
    variable r6271 : std_logic_vector(0 to 0) := (others => '0');
    variable r6270 : std_logic_vector(0 to 0) := (others => '0');
    variable r6269 : std_logic_vector(0 to 0) := (others => '0');
    variable r6268 : std_logic_vector(0 to 0) := (others => '0');
    variable r6267 : std_logic_vector(0 to 0) := (others => '0');
    variable r6266 : std_logic_vector(0 to 0) := (others => '0');
    variable r6265 : std_logic_vector(0 to 0) := (others => '0');
    variable r6264 : std_logic_vector(0 to 0) := (others => '0');
    variable r6263 : std_logic_vector(0 to 0) := (others => '0');
    variable r6262 : std_logic_vector(0 to 0) := (others => '0');
    variable r6261 : std_logic_vector(0 to 0) := (others => '0');
    variable r6260 : std_logic_vector(0 to 0) := (others => '0');
    variable r6259 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r6260 := "0";
    null;
    r6261 := (r6260);
    r6262 := "0";
    null;
    r6263 := (r6262);
    r6264 := "0";
    null;
    r6265 := (r6264);
    r6266 := "1";
    null;
    r6267 := (r6266);
    r6268 := "1";
    null;
    r6269 := (r6268);
    r6270 := "1";
    null;
    r6271 := (r6270);
    r6272 := "1";
    null;
    r6273 := (r6272);
    r6274 := "0";
    null;
    r6275 := (r6274);
    r6276 := "0";
    null;
    r6277 := (r6276);
    r6278 := "0";
    null;
    r6279 := (r6278);
    r6280 := "1";
    null;
    r6281 := (r6280);
    r6282 := "1";
    null;
    r6283 := (r6282);
    r6284 := "0";
    null;
    r6285 := (r6284);
    r6286 := "1";
    null;
    r6287 := (r6286);
    r6288 := "1";
    null;
    r6289 := (r6288);
    r6290 := "1";
    null;
    r6291 := (r6290);
    r6292 := "0";
    null;
    r6293 := (r6292);
    r6294 := "1";
    null;
    r6295 := (r6294);
    r6296 := "1";
    null;
    r6297 := (r6296);
    r6298 := "0";
    null;
    r6299 := (r6298);
    r6300 := "1";
    null;
    r6301 := (r6300);
    r6302 := "1";
    null;
    r6303 := (r6302);
    r6304 := "0";
    null;
    r6305 := (r6304);
    r6306 := "0";
    null;
    r6307 := (r6306);
    r6308 := "0";
    null;
    r6309 := (r6308);
    r6310 := "0";
    null;
    r6311 := (r6310);
    r6312 := "0";
    null;
    r6313 := (r6312);
    r6314 := "0";
    null;
    r6315 := (r6314);
    r6316 := "1";
    null;
    r6317 := (r6316);
    r6318 := "0";
    null;
    r6319 := (r6318);
    r6320 := "0";
    null;
    r6321 := (r6320);
    r6322 := "0";
    null;
    r6323 := (r6322);
    r6259 := (r6261 & r6263 & r6265 & r6267 & r6269 & r6271 & r6273 & r6275 & r6277 & r6279 & r6281 & r6283 & r6285 & r6287 & r6289 & r6291 & r6293 & r6295 & r6297 & r6299 & r6301 & r6303 & r6305 & r6307 & r6309 & r6311 & r6313 & r6315 & r6317 & r6319 & r6321 & r6323);
    return r6259;
  end rewire_MetaprogrammingRWw1e376c08_6258;
  function rewire_MetaprogrammingRWw19a4c116_6189 return std_logic_vector
  is
    variable r6254 : std_logic_vector(0 to 0) := (others => '0');
    variable r6253 : std_logic_vector(0 to 0) := (others => '0');
    variable r6252 : std_logic_vector(0 to 0) := (others => '0');
    variable r6251 : std_logic_vector(0 to 0) := (others => '0');
    variable r6250 : std_logic_vector(0 to 0) := (others => '0');
    variable r6249 : std_logic_vector(0 to 0) := (others => '0');
    variable r6248 : std_logic_vector(0 to 0) := (others => '0');
    variable r6247 : std_logic_vector(0 to 0) := (others => '0');
    variable r6246 : std_logic_vector(0 to 0) := (others => '0');
    variable r6245 : std_logic_vector(0 to 0) := (others => '0');
    variable r6244 : std_logic_vector(0 to 0) := (others => '0');
    variable r6243 : std_logic_vector(0 to 0) := (others => '0');
    variable r6242 : std_logic_vector(0 to 0) := (others => '0');
    variable r6241 : std_logic_vector(0 to 0) := (others => '0');
    variable r6240 : std_logic_vector(0 to 0) := (others => '0');
    variable r6239 : std_logic_vector(0 to 0) := (others => '0');
    variable r6238 : std_logic_vector(0 to 0) := (others => '0');
    variable r6237 : std_logic_vector(0 to 0) := (others => '0');
    variable r6236 : std_logic_vector(0 to 0) := (others => '0');
    variable r6235 : std_logic_vector(0 to 0) := (others => '0');
    variable r6234 : std_logic_vector(0 to 0) := (others => '0');
    variable r6233 : std_logic_vector(0 to 0) := (others => '0');
    variable r6232 : std_logic_vector(0 to 0) := (others => '0');
    variable r6231 : std_logic_vector(0 to 0) := (others => '0');
    variable r6230 : std_logic_vector(0 to 0) := (others => '0');
    variable r6229 : std_logic_vector(0 to 0) := (others => '0');
    variable r6228 : std_logic_vector(0 to 0) := (others => '0');
    variable r6227 : std_logic_vector(0 to 0) := (others => '0');
    variable r6226 : std_logic_vector(0 to 0) := (others => '0');
    variable r6225 : std_logic_vector(0 to 0) := (others => '0');
    variable r6224 : std_logic_vector(0 to 0) := (others => '0');
    variable r6223 : std_logic_vector(0 to 0) := (others => '0');
    variable r6222 : std_logic_vector(0 to 0) := (others => '0');
    variable r6221 : std_logic_vector(0 to 0) := (others => '0');
    variable r6220 : std_logic_vector(0 to 0) := (others => '0');
    variable r6219 : std_logic_vector(0 to 0) := (others => '0');
    variable r6218 : std_logic_vector(0 to 0) := (others => '0');
    variable r6217 : std_logic_vector(0 to 0) := (others => '0');
    variable r6216 : std_logic_vector(0 to 0) := (others => '0');
    variable r6215 : std_logic_vector(0 to 0) := (others => '0');
    variable r6214 : std_logic_vector(0 to 0) := (others => '0');
    variable r6213 : std_logic_vector(0 to 0) := (others => '0');
    variable r6212 : std_logic_vector(0 to 0) := (others => '0');
    variable r6211 : std_logic_vector(0 to 0) := (others => '0');
    variable r6210 : std_logic_vector(0 to 0) := (others => '0');
    variable r6209 : std_logic_vector(0 to 0) := (others => '0');
    variable r6208 : std_logic_vector(0 to 0) := (others => '0');
    variable r6207 : std_logic_vector(0 to 0) := (others => '0');
    variable r6206 : std_logic_vector(0 to 0) := (others => '0');
    variable r6205 : std_logic_vector(0 to 0) := (others => '0');
    variable r6204 : std_logic_vector(0 to 0) := (others => '0');
    variable r6203 : std_logic_vector(0 to 0) := (others => '0');
    variable r6202 : std_logic_vector(0 to 0) := (others => '0');
    variable r6201 : std_logic_vector(0 to 0) := (others => '0');
    variable r6200 : std_logic_vector(0 to 0) := (others => '0');
    variable r6199 : std_logic_vector(0 to 0) := (others => '0');
    variable r6198 : std_logic_vector(0 to 0) := (others => '0');
    variable r6197 : std_logic_vector(0 to 0) := (others => '0');
    variable r6196 : std_logic_vector(0 to 0) := (others => '0');
    variable r6195 : std_logic_vector(0 to 0) := (others => '0');
    variable r6194 : std_logic_vector(0 to 0) := (others => '0');
    variable r6193 : std_logic_vector(0 to 0) := (others => '0');
    variable r6192 : std_logic_vector(0 to 0) := (others => '0');
    variable r6191 : std_logic_vector(0 to 0) := (others => '0');
    variable r6190 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r6191 := "0";
    null;
    r6192 := (r6191);
    r6193 := "0";
    null;
    r6194 := (r6193);
    r6195 := "0";
    null;
    r6196 := (r6195);
    r6197 := "1";
    null;
    r6198 := (r6197);
    r6199 := "1";
    null;
    r6200 := (r6199);
    r6201 := "0";
    null;
    r6202 := (r6201);
    r6203 := "0";
    null;
    r6204 := (r6203);
    r6205 := "1";
    null;
    r6206 := (r6205);
    r6207 := "1";
    null;
    r6208 := (r6207);
    r6209 := "0";
    null;
    r6210 := (r6209);
    r6211 := "1";
    null;
    r6212 := (r6211);
    r6213 := "0";
    null;
    r6214 := (r6213);
    r6215 := "0";
    null;
    r6216 := (r6215);
    r6217 := "1";
    null;
    r6218 := (r6217);
    r6219 := "0";
    null;
    r6220 := (r6219);
    r6221 := "0";
    null;
    r6222 := (r6221);
    r6223 := "1";
    null;
    r6224 := (r6223);
    r6225 := "1";
    null;
    r6226 := (r6225);
    r6227 := "0";
    null;
    r6228 := (r6227);
    r6229 := "0";
    null;
    r6230 := (r6229);
    r6231 := "0";
    null;
    r6232 := (r6231);
    r6233 := "0";
    null;
    r6234 := (r6233);
    r6235 := "0";
    null;
    r6236 := (r6235);
    r6237 := "1";
    null;
    r6238 := (r6237);
    r6239 := "0";
    null;
    r6240 := (r6239);
    r6241 := "0";
    null;
    r6242 := (r6241);
    r6243 := "0";
    null;
    r6244 := (r6243);
    r6245 := "1";
    null;
    r6246 := (r6245);
    r6247 := "0";
    null;
    r6248 := (r6247);
    r6249 := "1";
    null;
    r6250 := (r6249);
    r6251 := "1";
    null;
    r6252 := (r6251);
    r6253 := "0";
    null;
    r6254 := (r6253);
    r6190 := (r6192 & r6194 & r6196 & r6198 & r6200 & r6202 & r6204 & r6206 & r6208 & r6210 & r6212 & r6214 & r6216 & r6218 & r6220 & r6222 & r6224 & r6226 & r6228 & r6230 & r6232 & r6234 & r6236 & r6238 & r6240 & r6242 & r6244 & r6246 & r6248 & r6250 & r6252 & r6254);
    return r6190;
  end rewire_MetaprogrammingRWw19a4c116_6189;
  function rewire_MetaprogrammingRWw106aa070_6120 return std_logic_vector
  is
    variable r6185 : std_logic_vector(0 to 0) := (others => '0');
    variable r6184 : std_logic_vector(0 to 0) := (others => '0');
    variable r6183 : std_logic_vector(0 to 0) := (others => '0');
    variable r6182 : std_logic_vector(0 to 0) := (others => '0');
    variable r6181 : std_logic_vector(0 to 0) := (others => '0');
    variable r6180 : std_logic_vector(0 to 0) := (others => '0');
    variable r6179 : std_logic_vector(0 to 0) := (others => '0');
    variable r6178 : std_logic_vector(0 to 0) := (others => '0');
    variable r6177 : std_logic_vector(0 to 0) := (others => '0');
    variable r6176 : std_logic_vector(0 to 0) := (others => '0');
    variable r6175 : std_logic_vector(0 to 0) := (others => '0');
    variable r6174 : std_logic_vector(0 to 0) := (others => '0');
    variable r6173 : std_logic_vector(0 to 0) := (others => '0');
    variable r6172 : std_logic_vector(0 to 0) := (others => '0');
    variable r6171 : std_logic_vector(0 to 0) := (others => '0');
    variable r6170 : std_logic_vector(0 to 0) := (others => '0');
    variable r6169 : std_logic_vector(0 to 0) := (others => '0');
    variable r6168 : std_logic_vector(0 to 0) := (others => '0');
    variable r6167 : std_logic_vector(0 to 0) := (others => '0');
    variable r6166 : std_logic_vector(0 to 0) := (others => '0');
    variable r6165 : std_logic_vector(0 to 0) := (others => '0');
    variable r6164 : std_logic_vector(0 to 0) := (others => '0');
    variable r6163 : std_logic_vector(0 to 0) := (others => '0');
    variable r6162 : std_logic_vector(0 to 0) := (others => '0');
    variable r6161 : std_logic_vector(0 to 0) := (others => '0');
    variable r6160 : std_logic_vector(0 to 0) := (others => '0');
    variable r6159 : std_logic_vector(0 to 0) := (others => '0');
    variable r6158 : std_logic_vector(0 to 0) := (others => '0');
    variable r6157 : std_logic_vector(0 to 0) := (others => '0');
    variable r6156 : std_logic_vector(0 to 0) := (others => '0');
    variable r6155 : std_logic_vector(0 to 0) := (others => '0');
    variable r6154 : std_logic_vector(0 to 0) := (others => '0');
    variable r6153 : std_logic_vector(0 to 0) := (others => '0');
    variable r6152 : std_logic_vector(0 to 0) := (others => '0');
    variable r6151 : std_logic_vector(0 to 0) := (others => '0');
    variable r6150 : std_logic_vector(0 to 0) := (others => '0');
    variable r6149 : std_logic_vector(0 to 0) := (others => '0');
    variable r6148 : std_logic_vector(0 to 0) := (others => '0');
    variable r6147 : std_logic_vector(0 to 0) := (others => '0');
    variable r6146 : std_logic_vector(0 to 0) := (others => '0');
    variable r6145 : std_logic_vector(0 to 0) := (others => '0');
    variable r6144 : std_logic_vector(0 to 0) := (others => '0');
    variable r6143 : std_logic_vector(0 to 0) := (others => '0');
    variable r6142 : std_logic_vector(0 to 0) := (others => '0');
    variable r6141 : std_logic_vector(0 to 0) := (others => '0');
    variable r6140 : std_logic_vector(0 to 0) := (others => '0');
    variable r6139 : std_logic_vector(0 to 0) := (others => '0');
    variable r6138 : std_logic_vector(0 to 0) := (others => '0');
    variable r6137 : std_logic_vector(0 to 0) := (others => '0');
    variable r6136 : std_logic_vector(0 to 0) := (others => '0');
    variable r6135 : std_logic_vector(0 to 0) := (others => '0');
    variable r6134 : std_logic_vector(0 to 0) := (others => '0');
    variable r6133 : std_logic_vector(0 to 0) := (others => '0');
    variable r6132 : std_logic_vector(0 to 0) := (others => '0');
    variable r6131 : std_logic_vector(0 to 0) := (others => '0');
    variable r6130 : std_logic_vector(0 to 0) := (others => '0');
    variable r6129 : std_logic_vector(0 to 0) := (others => '0');
    variable r6128 : std_logic_vector(0 to 0) := (others => '0');
    variable r6127 : std_logic_vector(0 to 0) := (others => '0');
    variable r6126 : std_logic_vector(0 to 0) := (others => '0');
    variable r6125 : std_logic_vector(0 to 0) := (others => '0');
    variable r6124 : std_logic_vector(0 to 0) := (others => '0');
    variable r6123 : std_logic_vector(0 to 0) := (others => '0');
    variable r6122 : std_logic_vector(0 to 0) := (others => '0');
    variable r6121 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r6122 := "0";
    null;
    r6123 := (r6122);
    r6124 := "0";
    null;
    r6125 := (r6124);
    r6126 := "0";
    null;
    r6127 := (r6126);
    r6128 := "1";
    null;
    r6129 := (r6128);
    r6130 := "0";
    null;
    r6131 := (r6130);
    r6132 := "0";
    null;
    r6133 := (r6132);
    r6134 := "0";
    null;
    r6135 := (r6134);
    r6136 := "0";
    null;
    r6137 := (r6136);
    r6138 := "0";
    null;
    r6139 := (r6138);
    r6140 := "1";
    null;
    r6141 := (r6140);
    r6142 := "1";
    null;
    r6143 := (r6142);
    r6144 := "0";
    null;
    r6145 := (r6144);
    r6146 := "1";
    null;
    r6147 := (r6146);
    r6148 := "0";
    null;
    r6149 := (r6148);
    r6150 := "1";
    null;
    r6151 := (r6150);
    r6152 := "0";
    null;
    r6153 := (r6152);
    r6154 := "1";
    null;
    r6155 := (r6154);
    r6156 := "0";
    null;
    r6157 := (r6156);
    r6158 := "1";
    null;
    r6159 := (r6158);
    r6160 := "0";
    null;
    r6161 := (r6160);
    r6162 := "0";
    null;
    r6163 := (r6162);
    r6164 := "0";
    null;
    r6165 := (r6164);
    r6166 := "0";
    null;
    r6167 := (r6166);
    r6168 := "0";
    null;
    r6169 := (r6168);
    r6170 := "0";
    null;
    r6171 := (r6170);
    r6172 := "1";
    null;
    r6173 := (r6172);
    r6174 := "1";
    null;
    r6175 := (r6174);
    r6176 := "1";
    null;
    r6177 := (r6176);
    r6178 := "0";
    null;
    r6179 := (r6178);
    r6180 := "0";
    null;
    r6181 := (r6180);
    r6182 := "0";
    null;
    r6183 := (r6182);
    r6184 := "0";
    null;
    r6185 := (r6184);
    r6121 := (r6123 & r6125 & r6127 & r6129 & r6131 & r6133 & r6135 & r6137 & r6139 & r6141 & r6143 & r6145 & r6147 & r6149 & r6151 & r6153 & r6155 & r6157 & r6159 & r6161 & r6163 & r6165 & r6167 & r6169 & r6171 & r6173 & r6175 & r6177 & r6179 & r6181 & r6183 & r6185);
    return r6121;
  end rewire_MetaprogrammingRWw106aa070_6120;
  function rewire_MetaprogrammingRWwf40e3585_6051 return std_logic_vector
  is
    variable r6116 : std_logic_vector(0 to 0) := (others => '0');
    variable r6115 : std_logic_vector(0 to 0) := (others => '0');
    variable r6114 : std_logic_vector(0 to 0) := (others => '0');
    variable r6113 : std_logic_vector(0 to 0) := (others => '0');
    variable r6112 : std_logic_vector(0 to 0) := (others => '0');
    variable r6111 : std_logic_vector(0 to 0) := (others => '0');
    variable r6110 : std_logic_vector(0 to 0) := (others => '0');
    variable r6109 : std_logic_vector(0 to 0) := (others => '0');
    variable r6108 : std_logic_vector(0 to 0) := (others => '0');
    variable r6107 : std_logic_vector(0 to 0) := (others => '0');
    variable r6106 : std_logic_vector(0 to 0) := (others => '0');
    variable r6105 : std_logic_vector(0 to 0) := (others => '0');
    variable r6104 : std_logic_vector(0 to 0) := (others => '0');
    variable r6103 : std_logic_vector(0 to 0) := (others => '0');
    variable r6102 : std_logic_vector(0 to 0) := (others => '0');
    variable r6101 : std_logic_vector(0 to 0) := (others => '0');
    variable r6100 : std_logic_vector(0 to 0) := (others => '0');
    variable r6099 : std_logic_vector(0 to 0) := (others => '0');
    variable r6098 : std_logic_vector(0 to 0) := (others => '0');
    variable r6097 : std_logic_vector(0 to 0) := (others => '0');
    variable r6096 : std_logic_vector(0 to 0) := (others => '0');
    variable r6095 : std_logic_vector(0 to 0) := (others => '0');
    variable r6094 : std_logic_vector(0 to 0) := (others => '0');
    variable r6093 : std_logic_vector(0 to 0) := (others => '0');
    variable r6092 : std_logic_vector(0 to 0) := (others => '0');
    variable r6091 : std_logic_vector(0 to 0) := (others => '0');
    variable r6090 : std_logic_vector(0 to 0) := (others => '0');
    variable r6089 : std_logic_vector(0 to 0) := (others => '0');
    variable r6088 : std_logic_vector(0 to 0) := (others => '0');
    variable r6087 : std_logic_vector(0 to 0) := (others => '0');
    variable r6086 : std_logic_vector(0 to 0) := (others => '0');
    variable r6085 : std_logic_vector(0 to 0) := (others => '0');
    variable r6084 : std_logic_vector(0 to 0) := (others => '0');
    variable r6083 : std_logic_vector(0 to 0) := (others => '0');
    variable r6082 : std_logic_vector(0 to 0) := (others => '0');
    variable r6081 : std_logic_vector(0 to 0) := (others => '0');
    variable r6080 : std_logic_vector(0 to 0) := (others => '0');
    variable r6079 : std_logic_vector(0 to 0) := (others => '0');
    variable r6078 : std_logic_vector(0 to 0) := (others => '0');
    variable r6077 : std_logic_vector(0 to 0) := (others => '0');
    variable r6076 : std_logic_vector(0 to 0) := (others => '0');
    variable r6075 : std_logic_vector(0 to 0) := (others => '0');
    variable r6074 : std_logic_vector(0 to 0) := (others => '0');
    variable r6073 : std_logic_vector(0 to 0) := (others => '0');
    variable r6072 : std_logic_vector(0 to 0) := (others => '0');
    variable r6071 : std_logic_vector(0 to 0) := (others => '0');
    variable r6070 : std_logic_vector(0 to 0) := (others => '0');
    variable r6069 : std_logic_vector(0 to 0) := (others => '0');
    variable r6068 : std_logic_vector(0 to 0) := (others => '0');
    variable r6067 : std_logic_vector(0 to 0) := (others => '0');
    variable r6066 : std_logic_vector(0 to 0) := (others => '0');
    variable r6065 : std_logic_vector(0 to 0) := (others => '0');
    variable r6064 : std_logic_vector(0 to 0) := (others => '0');
    variable r6063 : std_logic_vector(0 to 0) := (others => '0');
    variable r6062 : std_logic_vector(0 to 0) := (others => '0');
    variable r6061 : std_logic_vector(0 to 0) := (others => '0');
    variable r6060 : std_logic_vector(0 to 0) := (others => '0');
    variable r6059 : std_logic_vector(0 to 0) := (others => '0');
    variable r6058 : std_logic_vector(0 to 0) := (others => '0');
    variable r6057 : std_logic_vector(0 to 0) := (others => '0');
    variable r6056 : std_logic_vector(0 to 0) := (others => '0');
    variable r6055 : std_logic_vector(0 to 0) := (others => '0');
    variable r6054 : std_logic_vector(0 to 0) := (others => '0');
    variable r6053 : std_logic_vector(0 to 0) := (others => '0');
    variable r6052 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r6053 := "1";
    null;
    r6054 := (r6053);
    r6055 := "1";
    null;
    r6056 := (r6055);
    r6057 := "1";
    null;
    r6058 := (r6057);
    r6059 := "1";
    null;
    r6060 := (r6059);
    r6061 := "0";
    null;
    r6062 := (r6061);
    r6063 := "1";
    null;
    r6064 := (r6063);
    r6065 := "0";
    null;
    r6066 := (r6065);
    r6067 := "0";
    null;
    r6068 := (r6067);
    r6069 := "0";
    null;
    r6070 := (r6069);
    r6071 := "0";
    null;
    r6072 := (r6071);
    r6073 := "0";
    null;
    r6074 := (r6073);
    r6075 := "0";
    null;
    r6076 := (r6075);
    r6077 := "1";
    null;
    r6078 := (r6077);
    r6079 := "1";
    null;
    r6080 := (r6079);
    r6081 := "1";
    null;
    r6082 := (r6081);
    r6083 := "0";
    null;
    r6084 := (r6083);
    r6085 := "0";
    null;
    r6086 := (r6085);
    r6087 := "0";
    null;
    r6088 := (r6087);
    r6089 := "1";
    null;
    r6090 := (r6089);
    r6091 := "1";
    null;
    r6092 := (r6091);
    r6093 := "0";
    null;
    r6094 := (r6093);
    r6095 := "1";
    null;
    r6096 := (r6095);
    r6097 := "0";
    null;
    r6098 := (r6097);
    r6099 := "1";
    null;
    r6100 := (r6099);
    r6101 := "1";
    null;
    r6102 := (r6101);
    r6103 := "0";
    null;
    r6104 := (r6103);
    r6105 := "0";
    null;
    r6106 := (r6105);
    r6107 := "0";
    null;
    r6108 := (r6107);
    r6109 := "0";
    null;
    r6110 := (r6109);
    r6111 := "1";
    null;
    r6112 := (r6111);
    r6113 := "0";
    null;
    r6114 := (r6113);
    r6115 := "1";
    null;
    r6116 := (r6115);
    r6052 := (r6054 & r6056 & r6058 & r6060 & r6062 & r6064 & r6066 & r6068 & r6070 & r6072 & r6074 & r6076 & r6078 & r6080 & r6082 & r6084 & r6086 & r6088 & r6090 & r6092 & r6094 & r6096 & r6098 & r6100 & r6102 & r6104 & r6106 & r6108 & r6110 & r6112 & r6114 & r6116);
    return r6052;
  end rewire_MetaprogrammingRWwf40e3585_6051;
  function rewire_MetaprogrammingRWwd6990624_5982 return std_logic_vector
  is
    variable r6047 : std_logic_vector(0 to 0) := (others => '0');
    variable r6046 : std_logic_vector(0 to 0) := (others => '0');
    variable r6045 : std_logic_vector(0 to 0) := (others => '0');
    variable r6044 : std_logic_vector(0 to 0) := (others => '0');
    variable r6043 : std_logic_vector(0 to 0) := (others => '0');
    variable r6042 : std_logic_vector(0 to 0) := (others => '0');
    variable r6041 : std_logic_vector(0 to 0) := (others => '0');
    variable r6040 : std_logic_vector(0 to 0) := (others => '0');
    variable r6039 : std_logic_vector(0 to 0) := (others => '0');
    variable r6038 : std_logic_vector(0 to 0) := (others => '0');
    variable r6037 : std_logic_vector(0 to 0) := (others => '0');
    variable r6036 : std_logic_vector(0 to 0) := (others => '0');
    variable r6035 : std_logic_vector(0 to 0) := (others => '0');
    variable r6034 : std_logic_vector(0 to 0) := (others => '0');
    variable r6033 : std_logic_vector(0 to 0) := (others => '0');
    variable r6032 : std_logic_vector(0 to 0) := (others => '0');
    variable r6031 : std_logic_vector(0 to 0) := (others => '0');
    variable r6030 : std_logic_vector(0 to 0) := (others => '0');
    variable r6029 : std_logic_vector(0 to 0) := (others => '0');
    variable r6028 : std_logic_vector(0 to 0) := (others => '0');
    variable r6027 : std_logic_vector(0 to 0) := (others => '0');
    variable r6026 : std_logic_vector(0 to 0) := (others => '0');
    variable r6025 : std_logic_vector(0 to 0) := (others => '0');
    variable r6024 : std_logic_vector(0 to 0) := (others => '0');
    variable r6023 : std_logic_vector(0 to 0) := (others => '0');
    variable r6022 : std_logic_vector(0 to 0) := (others => '0');
    variable r6021 : std_logic_vector(0 to 0) := (others => '0');
    variable r6020 : std_logic_vector(0 to 0) := (others => '0');
    variable r6019 : std_logic_vector(0 to 0) := (others => '0');
    variable r6018 : std_logic_vector(0 to 0) := (others => '0');
    variable r6017 : std_logic_vector(0 to 0) := (others => '0');
    variable r6016 : std_logic_vector(0 to 0) := (others => '0');
    variable r6015 : std_logic_vector(0 to 0) := (others => '0');
    variable r6014 : std_logic_vector(0 to 0) := (others => '0');
    variable r6013 : std_logic_vector(0 to 0) := (others => '0');
    variable r6012 : std_logic_vector(0 to 0) := (others => '0');
    variable r6011 : std_logic_vector(0 to 0) := (others => '0');
    variable r6010 : std_logic_vector(0 to 0) := (others => '0');
    variable r6009 : std_logic_vector(0 to 0) := (others => '0');
    variable r6008 : std_logic_vector(0 to 0) := (others => '0');
    variable r6007 : std_logic_vector(0 to 0) := (others => '0');
    variable r6006 : std_logic_vector(0 to 0) := (others => '0');
    variable r6005 : std_logic_vector(0 to 0) := (others => '0');
    variable r6004 : std_logic_vector(0 to 0) := (others => '0');
    variable r6003 : std_logic_vector(0 to 0) := (others => '0');
    variable r6002 : std_logic_vector(0 to 0) := (others => '0');
    variable r6001 : std_logic_vector(0 to 0) := (others => '0');
    variable r6000 : std_logic_vector(0 to 0) := (others => '0');
    variable r5999 : std_logic_vector(0 to 0) := (others => '0');
    variable r5998 : std_logic_vector(0 to 0) := (others => '0');
    variable r5997 : std_logic_vector(0 to 0) := (others => '0');
    variable r5996 : std_logic_vector(0 to 0) := (others => '0');
    variable r5995 : std_logic_vector(0 to 0) := (others => '0');
    variable r5994 : std_logic_vector(0 to 0) := (others => '0');
    variable r5993 : std_logic_vector(0 to 0) := (others => '0');
    variable r5992 : std_logic_vector(0 to 0) := (others => '0');
    variable r5991 : std_logic_vector(0 to 0) := (others => '0');
    variable r5990 : std_logic_vector(0 to 0) := (others => '0');
    variable r5989 : std_logic_vector(0 to 0) := (others => '0');
    variable r5988 : std_logic_vector(0 to 0) := (others => '0');
    variable r5987 : std_logic_vector(0 to 0) := (others => '0');
    variable r5986 : std_logic_vector(0 to 0) := (others => '0');
    variable r5985 : std_logic_vector(0 to 0) := (others => '0');
    variable r5984 : std_logic_vector(0 to 0) := (others => '0');
    variable r5983 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r5984 := "1";
    null;
    r5985 := (r5984);
    r5986 := "1";
    null;
    r5987 := (r5986);
    r5988 := "0";
    null;
    r5989 := (r5988);
    r5990 := "1";
    null;
    r5991 := (r5990);
    r5992 := "0";
    null;
    r5993 := (r5992);
    r5994 := "1";
    null;
    r5995 := (r5994);
    r5996 := "1";
    null;
    r5997 := (r5996);
    r5998 := "0";
    null;
    r5999 := (r5998);
    r6000 := "1";
    null;
    r6001 := (r6000);
    r6002 := "0";
    null;
    r6003 := (r6002);
    r6004 := "0";
    null;
    r6005 := (r6004);
    r6006 := "1";
    null;
    r6007 := (r6006);
    r6008 := "1";
    null;
    r6009 := (r6008);
    r6010 := "0";
    null;
    r6011 := (r6010);
    r6012 := "0";
    null;
    r6013 := (r6012);
    r6014 := "1";
    null;
    r6015 := (r6014);
    r6016 := "0";
    null;
    r6017 := (r6016);
    r6018 := "0";
    null;
    r6019 := (r6018);
    r6020 := "0";
    null;
    r6021 := (r6020);
    r6022 := "0";
    null;
    r6023 := (r6022);
    r6024 := "0";
    null;
    r6025 := (r6024);
    r6026 := "1";
    null;
    r6027 := (r6026);
    r6028 := "1";
    null;
    r6029 := (r6028);
    r6030 := "0";
    null;
    r6031 := (r6030);
    r6032 := "0";
    null;
    r6033 := (r6032);
    r6034 := "0";
    null;
    r6035 := (r6034);
    r6036 := "1";
    null;
    r6037 := (r6036);
    r6038 := "0";
    null;
    r6039 := (r6038);
    r6040 := "0";
    null;
    r6041 := (r6040);
    r6042 := "1";
    null;
    r6043 := (r6042);
    r6044 := "0";
    null;
    r6045 := (r6044);
    r6046 := "0";
    null;
    r6047 := (r6046);
    r5983 := (r5985 & r5987 & r5989 & r5991 & r5993 & r5995 & r5997 & r5999 & r6001 & r6003 & r6005 & r6007 & r6009 & r6011 & r6013 & r6015 & r6017 & r6019 & r6021 & r6023 & r6025 & r6027 & r6029 & r6031 & r6033 & r6035 & r6037 & r6039 & r6041 & r6043 & r6045 & r6047);
    return r5983;
  end rewire_MetaprogrammingRWwd6990624_5982;
  function rewire_MetaprogrammingRWwd192e819_5913 return std_logic_vector
  is
    variable r5978 : std_logic_vector(0 to 0) := (others => '0');
    variable r5977 : std_logic_vector(0 to 0) := (others => '0');
    variable r5976 : std_logic_vector(0 to 0) := (others => '0');
    variable r5975 : std_logic_vector(0 to 0) := (others => '0');
    variable r5974 : std_logic_vector(0 to 0) := (others => '0');
    variable r5973 : std_logic_vector(0 to 0) := (others => '0');
    variable r5972 : std_logic_vector(0 to 0) := (others => '0');
    variable r5971 : std_logic_vector(0 to 0) := (others => '0');
    variable r5970 : std_logic_vector(0 to 0) := (others => '0');
    variable r5969 : std_logic_vector(0 to 0) := (others => '0');
    variable r5968 : std_logic_vector(0 to 0) := (others => '0');
    variable r5967 : std_logic_vector(0 to 0) := (others => '0');
    variable r5966 : std_logic_vector(0 to 0) := (others => '0');
    variable r5965 : std_logic_vector(0 to 0) := (others => '0');
    variable r5964 : std_logic_vector(0 to 0) := (others => '0');
    variable r5963 : std_logic_vector(0 to 0) := (others => '0');
    variable r5962 : std_logic_vector(0 to 0) := (others => '0');
    variable r5961 : std_logic_vector(0 to 0) := (others => '0');
    variable r5960 : std_logic_vector(0 to 0) := (others => '0');
    variable r5959 : std_logic_vector(0 to 0) := (others => '0');
    variable r5958 : std_logic_vector(0 to 0) := (others => '0');
    variable r5957 : std_logic_vector(0 to 0) := (others => '0');
    variable r5956 : std_logic_vector(0 to 0) := (others => '0');
    variable r5955 : std_logic_vector(0 to 0) := (others => '0');
    variable r5954 : std_logic_vector(0 to 0) := (others => '0');
    variable r5953 : std_logic_vector(0 to 0) := (others => '0');
    variable r5952 : std_logic_vector(0 to 0) := (others => '0');
    variable r5951 : std_logic_vector(0 to 0) := (others => '0');
    variable r5950 : std_logic_vector(0 to 0) := (others => '0');
    variable r5949 : std_logic_vector(0 to 0) := (others => '0');
    variable r5948 : std_logic_vector(0 to 0) := (others => '0');
    variable r5947 : std_logic_vector(0 to 0) := (others => '0');
    variable r5946 : std_logic_vector(0 to 0) := (others => '0');
    variable r5945 : std_logic_vector(0 to 0) := (others => '0');
    variable r5944 : std_logic_vector(0 to 0) := (others => '0');
    variable r5943 : std_logic_vector(0 to 0) := (others => '0');
    variable r5942 : std_logic_vector(0 to 0) := (others => '0');
    variable r5941 : std_logic_vector(0 to 0) := (others => '0');
    variable r5940 : std_logic_vector(0 to 0) := (others => '0');
    variable r5939 : std_logic_vector(0 to 0) := (others => '0');
    variable r5938 : std_logic_vector(0 to 0) := (others => '0');
    variable r5937 : std_logic_vector(0 to 0) := (others => '0');
    variable r5936 : std_logic_vector(0 to 0) := (others => '0');
    variable r5935 : std_logic_vector(0 to 0) := (others => '0');
    variable r5934 : std_logic_vector(0 to 0) := (others => '0');
    variable r5933 : std_logic_vector(0 to 0) := (others => '0');
    variable r5932 : std_logic_vector(0 to 0) := (others => '0');
    variable r5931 : std_logic_vector(0 to 0) := (others => '0');
    variable r5930 : std_logic_vector(0 to 0) := (others => '0');
    variable r5929 : std_logic_vector(0 to 0) := (others => '0');
    variable r5928 : std_logic_vector(0 to 0) := (others => '0');
    variable r5927 : std_logic_vector(0 to 0) := (others => '0');
    variable r5926 : std_logic_vector(0 to 0) := (others => '0');
    variable r5925 : std_logic_vector(0 to 0) := (others => '0');
    variable r5924 : std_logic_vector(0 to 0) := (others => '0');
    variable r5923 : std_logic_vector(0 to 0) := (others => '0');
    variable r5922 : std_logic_vector(0 to 0) := (others => '0');
    variable r5921 : std_logic_vector(0 to 0) := (others => '0');
    variable r5920 : std_logic_vector(0 to 0) := (others => '0');
    variable r5919 : std_logic_vector(0 to 0) := (others => '0');
    variable r5918 : std_logic_vector(0 to 0) := (others => '0');
    variable r5917 : std_logic_vector(0 to 0) := (others => '0');
    variable r5916 : std_logic_vector(0 to 0) := (others => '0');
    variable r5915 : std_logic_vector(0 to 0) := (others => '0');
    variable r5914 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r5915 := "1";
    null;
    r5916 := (r5915);
    r5917 := "1";
    null;
    r5918 := (r5917);
    r5919 := "0";
    null;
    r5920 := (r5919);
    r5921 := "1";
    null;
    r5922 := (r5921);
    r5923 := "0";
    null;
    r5924 := (r5923);
    r5925 := "0";
    null;
    r5926 := (r5925);
    r5927 := "0";
    null;
    r5928 := (r5927);
    r5929 := "1";
    null;
    r5930 := (r5929);
    r5931 := "1";
    null;
    r5932 := (r5931);
    r5933 := "0";
    null;
    r5934 := (r5933);
    r5935 := "0";
    null;
    r5936 := (r5935);
    r5937 := "1";
    null;
    r5938 := (r5937);
    r5939 := "0";
    null;
    r5940 := (r5939);
    r5941 := "0";
    null;
    r5942 := (r5941);
    r5943 := "1";
    null;
    r5944 := (r5943);
    r5945 := "0";
    null;
    r5946 := (r5945);
    r5947 := "1";
    null;
    r5948 := (r5947);
    r5949 := "1";
    null;
    r5950 := (r5949);
    r5951 := "1";
    null;
    r5952 := (r5951);
    r5953 := "0";
    null;
    r5954 := (r5953);
    r5955 := "1";
    null;
    r5956 := (r5955);
    r5957 := "0";
    null;
    r5958 := (r5957);
    r5959 := "0";
    null;
    r5960 := (r5959);
    r5961 := "0";
    null;
    r5962 := (r5961);
    r5963 := "0";
    null;
    r5964 := (r5963);
    r5965 := "0";
    null;
    r5966 := (r5965);
    r5967 := "0";
    null;
    r5968 := (r5967);
    r5969 := "1";
    null;
    r5970 := (r5969);
    r5971 := "1";
    null;
    r5972 := (r5971);
    r5973 := "0";
    null;
    r5974 := (r5973);
    r5975 := "0";
    null;
    r5976 := (r5975);
    r5977 := "1";
    null;
    r5978 := (r5977);
    r5914 := (r5916 & r5918 & r5920 & r5922 & r5924 & r5926 & r5928 & r5930 & r5932 & r5934 & r5936 & r5938 & r5940 & r5942 & r5944 & r5946 & r5948 & r5950 & r5952 & r5954 & r5956 & r5958 & r5960 & r5962 & r5964 & r5966 & r5968 & r5970 & r5972 & r5974 & r5976 & r5978);
    return r5914;
  end rewire_MetaprogrammingRWwd192e819_5913;
  function rewire_MetaprogrammingRWwc76c51a3_5844 return std_logic_vector
  is
    variable r5909 : std_logic_vector(0 to 0) := (others => '0');
    variable r5908 : std_logic_vector(0 to 0) := (others => '0');
    variable r5907 : std_logic_vector(0 to 0) := (others => '0');
    variable r5906 : std_logic_vector(0 to 0) := (others => '0');
    variable r5905 : std_logic_vector(0 to 0) := (others => '0');
    variable r5904 : std_logic_vector(0 to 0) := (others => '0');
    variable r5903 : std_logic_vector(0 to 0) := (others => '0');
    variable r5902 : std_logic_vector(0 to 0) := (others => '0');
    variable r5901 : std_logic_vector(0 to 0) := (others => '0');
    variable r5900 : std_logic_vector(0 to 0) := (others => '0');
    variable r5899 : std_logic_vector(0 to 0) := (others => '0');
    variable r5898 : std_logic_vector(0 to 0) := (others => '0');
    variable r5897 : std_logic_vector(0 to 0) := (others => '0');
    variable r5896 : std_logic_vector(0 to 0) := (others => '0');
    variable r5895 : std_logic_vector(0 to 0) := (others => '0');
    variable r5894 : std_logic_vector(0 to 0) := (others => '0');
    variable r5893 : std_logic_vector(0 to 0) := (others => '0');
    variable r5892 : std_logic_vector(0 to 0) := (others => '0');
    variable r5891 : std_logic_vector(0 to 0) := (others => '0');
    variable r5890 : std_logic_vector(0 to 0) := (others => '0');
    variable r5889 : std_logic_vector(0 to 0) := (others => '0');
    variable r5888 : std_logic_vector(0 to 0) := (others => '0');
    variable r5887 : std_logic_vector(0 to 0) := (others => '0');
    variable r5886 : std_logic_vector(0 to 0) := (others => '0');
    variable r5885 : std_logic_vector(0 to 0) := (others => '0');
    variable r5884 : std_logic_vector(0 to 0) := (others => '0');
    variable r5883 : std_logic_vector(0 to 0) := (others => '0');
    variable r5882 : std_logic_vector(0 to 0) := (others => '0');
    variable r5881 : std_logic_vector(0 to 0) := (others => '0');
    variable r5880 : std_logic_vector(0 to 0) := (others => '0');
    variable r5879 : std_logic_vector(0 to 0) := (others => '0');
    variable r5878 : std_logic_vector(0 to 0) := (others => '0');
    variable r5877 : std_logic_vector(0 to 0) := (others => '0');
    variable r5876 : std_logic_vector(0 to 0) := (others => '0');
    variable r5875 : std_logic_vector(0 to 0) := (others => '0');
    variable r5874 : std_logic_vector(0 to 0) := (others => '0');
    variable r5873 : std_logic_vector(0 to 0) := (others => '0');
    variable r5872 : std_logic_vector(0 to 0) := (others => '0');
    variable r5871 : std_logic_vector(0 to 0) := (others => '0');
    variable r5870 : std_logic_vector(0 to 0) := (others => '0');
    variable r5869 : std_logic_vector(0 to 0) := (others => '0');
    variable r5868 : std_logic_vector(0 to 0) := (others => '0');
    variable r5867 : std_logic_vector(0 to 0) := (others => '0');
    variable r5866 : std_logic_vector(0 to 0) := (others => '0');
    variable r5865 : std_logic_vector(0 to 0) := (others => '0');
    variable r5864 : std_logic_vector(0 to 0) := (others => '0');
    variable r5863 : std_logic_vector(0 to 0) := (others => '0');
    variable r5862 : std_logic_vector(0 to 0) := (others => '0');
    variable r5861 : std_logic_vector(0 to 0) := (others => '0');
    variable r5860 : std_logic_vector(0 to 0) := (others => '0');
    variable r5859 : std_logic_vector(0 to 0) := (others => '0');
    variable r5858 : std_logic_vector(0 to 0) := (others => '0');
    variable r5857 : std_logic_vector(0 to 0) := (others => '0');
    variable r5856 : std_logic_vector(0 to 0) := (others => '0');
    variable r5855 : std_logic_vector(0 to 0) := (others => '0');
    variable r5854 : std_logic_vector(0 to 0) := (others => '0');
    variable r5853 : std_logic_vector(0 to 0) := (others => '0');
    variable r5852 : std_logic_vector(0 to 0) := (others => '0');
    variable r5851 : std_logic_vector(0 to 0) := (others => '0');
    variable r5850 : std_logic_vector(0 to 0) := (others => '0');
    variable r5849 : std_logic_vector(0 to 0) := (others => '0');
    variable r5848 : std_logic_vector(0 to 0) := (others => '0');
    variable r5847 : std_logic_vector(0 to 0) := (others => '0');
    variable r5846 : std_logic_vector(0 to 0) := (others => '0');
    variable r5845 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r5846 := "1";
    null;
    r5847 := (r5846);
    r5848 := "1";
    null;
    r5849 := (r5848);
    r5850 := "0";
    null;
    r5851 := (r5850);
    r5852 := "0";
    null;
    r5853 := (r5852);
    r5854 := "0";
    null;
    r5855 := (r5854);
    r5856 := "1";
    null;
    r5857 := (r5856);
    r5858 := "1";
    null;
    r5859 := (r5858);
    r5860 := "1";
    null;
    r5861 := (r5860);
    r5862 := "0";
    null;
    r5863 := (r5862);
    r5864 := "1";
    null;
    r5865 := (r5864);
    r5866 := "1";
    null;
    r5867 := (r5866);
    r5868 := "0";
    null;
    r5869 := (r5868);
    r5870 := "1";
    null;
    r5871 := (r5870);
    r5872 := "1";
    null;
    r5873 := (r5872);
    r5874 := "0";
    null;
    r5875 := (r5874);
    r5876 := "0";
    null;
    r5877 := (r5876);
    r5878 := "0";
    null;
    r5879 := (r5878);
    r5880 := "1";
    null;
    r5881 := (r5880);
    r5882 := "0";
    null;
    r5883 := (r5882);
    r5884 := "1";
    null;
    r5885 := (r5884);
    r5886 := "0";
    null;
    r5887 := (r5886);
    r5888 := "0";
    null;
    r5889 := (r5888);
    r5890 := "0";
    null;
    r5891 := (r5890);
    r5892 := "1";
    null;
    r5893 := (r5892);
    r5894 := "1";
    null;
    r5895 := (r5894);
    r5896 := "0";
    null;
    r5897 := (r5896);
    r5898 := "1";
    null;
    r5899 := (r5898);
    r5900 := "0";
    null;
    r5901 := (r5900);
    r5902 := "0";
    null;
    r5903 := (r5902);
    r5904 := "0";
    null;
    r5905 := (r5904);
    r5906 := "1";
    null;
    r5907 := (r5906);
    r5908 := "1";
    null;
    r5909 := (r5908);
    r5845 := (r5847 & r5849 & r5851 & r5853 & r5855 & r5857 & r5859 & r5861 & r5863 & r5865 & r5867 & r5869 & r5871 & r5873 & r5875 & r5877 & r5879 & r5881 & r5883 & r5885 & r5887 & r5889 & r5891 & r5893 & r5895 & r5897 & r5899 & r5901 & r5903 & r5905 & r5907 & r5909);
    return r5845;
  end rewire_MetaprogrammingRWwc76c51a3_5844;
  function rewire_MetaprogrammingRWwc24b8b70_5775 return std_logic_vector
  is
    variable r5840 : std_logic_vector(0 to 0) := (others => '0');
    variable r5839 : std_logic_vector(0 to 0) := (others => '0');
    variable r5838 : std_logic_vector(0 to 0) := (others => '0');
    variable r5837 : std_logic_vector(0 to 0) := (others => '0');
    variable r5836 : std_logic_vector(0 to 0) := (others => '0');
    variable r5835 : std_logic_vector(0 to 0) := (others => '0');
    variable r5834 : std_logic_vector(0 to 0) := (others => '0');
    variable r5833 : std_logic_vector(0 to 0) := (others => '0');
    variable r5832 : std_logic_vector(0 to 0) := (others => '0');
    variable r5831 : std_logic_vector(0 to 0) := (others => '0');
    variable r5830 : std_logic_vector(0 to 0) := (others => '0');
    variable r5829 : std_logic_vector(0 to 0) := (others => '0');
    variable r5828 : std_logic_vector(0 to 0) := (others => '0');
    variable r5827 : std_logic_vector(0 to 0) := (others => '0');
    variable r5826 : std_logic_vector(0 to 0) := (others => '0');
    variable r5825 : std_logic_vector(0 to 0) := (others => '0');
    variable r5824 : std_logic_vector(0 to 0) := (others => '0');
    variable r5823 : std_logic_vector(0 to 0) := (others => '0');
    variable r5822 : std_logic_vector(0 to 0) := (others => '0');
    variable r5821 : std_logic_vector(0 to 0) := (others => '0');
    variable r5820 : std_logic_vector(0 to 0) := (others => '0');
    variable r5819 : std_logic_vector(0 to 0) := (others => '0');
    variable r5818 : std_logic_vector(0 to 0) := (others => '0');
    variable r5817 : std_logic_vector(0 to 0) := (others => '0');
    variable r5816 : std_logic_vector(0 to 0) := (others => '0');
    variable r5815 : std_logic_vector(0 to 0) := (others => '0');
    variable r5814 : std_logic_vector(0 to 0) := (others => '0');
    variable r5813 : std_logic_vector(0 to 0) := (others => '0');
    variable r5812 : std_logic_vector(0 to 0) := (others => '0');
    variable r5811 : std_logic_vector(0 to 0) := (others => '0');
    variable r5810 : std_logic_vector(0 to 0) := (others => '0');
    variable r5809 : std_logic_vector(0 to 0) := (others => '0');
    variable r5808 : std_logic_vector(0 to 0) := (others => '0');
    variable r5807 : std_logic_vector(0 to 0) := (others => '0');
    variable r5806 : std_logic_vector(0 to 0) := (others => '0');
    variable r5805 : std_logic_vector(0 to 0) := (others => '0');
    variable r5804 : std_logic_vector(0 to 0) := (others => '0');
    variable r5803 : std_logic_vector(0 to 0) := (others => '0');
    variable r5802 : std_logic_vector(0 to 0) := (others => '0');
    variable r5801 : std_logic_vector(0 to 0) := (others => '0');
    variable r5800 : std_logic_vector(0 to 0) := (others => '0');
    variable r5799 : std_logic_vector(0 to 0) := (others => '0');
    variable r5798 : std_logic_vector(0 to 0) := (others => '0');
    variable r5797 : std_logic_vector(0 to 0) := (others => '0');
    variable r5796 : std_logic_vector(0 to 0) := (others => '0');
    variable r5795 : std_logic_vector(0 to 0) := (others => '0');
    variable r5794 : std_logic_vector(0 to 0) := (others => '0');
    variable r5793 : std_logic_vector(0 to 0) := (others => '0');
    variable r5792 : std_logic_vector(0 to 0) := (others => '0');
    variable r5791 : std_logic_vector(0 to 0) := (others => '0');
    variable r5790 : std_logic_vector(0 to 0) := (others => '0');
    variable r5789 : std_logic_vector(0 to 0) := (others => '0');
    variable r5788 : std_logic_vector(0 to 0) := (others => '0');
    variable r5787 : std_logic_vector(0 to 0) := (others => '0');
    variable r5786 : std_logic_vector(0 to 0) := (others => '0');
    variable r5785 : std_logic_vector(0 to 0) := (others => '0');
    variable r5784 : std_logic_vector(0 to 0) := (others => '0');
    variable r5783 : std_logic_vector(0 to 0) := (others => '0');
    variable r5782 : std_logic_vector(0 to 0) := (others => '0');
    variable r5781 : std_logic_vector(0 to 0) := (others => '0');
    variable r5780 : std_logic_vector(0 to 0) := (others => '0');
    variable r5779 : std_logic_vector(0 to 0) := (others => '0');
    variable r5778 : std_logic_vector(0 to 0) := (others => '0');
    variable r5777 : std_logic_vector(0 to 0) := (others => '0');
    variable r5776 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r5777 := "1";
    null;
    r5778 := (r5777);
    r5779 := "1";
    null;
    r5780 := (r5779);
    r5781 := "0";
    null;
    r5782 := (r5781);
    r5783 := "0";
    null;
    r5784 := (r5783);
    r5785 := "0";
    null;
    r5786 := (r5785);
    r5787 := "0";
    null;
    r5788 := (r5787);
    r5789 := "1";
    null;
    r5790 := (r5789);
    r5791 := "0";
    null;
    r5792 := (r5791);
    r5793 := "0";
    null;
    r5794 := (r5793);
    r5795 := "1";
    null;
    r5796 := (r5795);
    r5797 := "0";
    null;
    r5798 := (r5797);
    r5799 := "0";
    null;
    r5800 := (r5799);
    r5801 := "1";
    null;
    r5802 := (r5801);
    r5803 := "0";
    null;
    r5804 := (r5803);
    r5805 := "1";
    null;
    r5806 := (r5805);
    r5807 := "1";
    null;
    r5808 := (r5807);
    r5809 := "1";
    null;
    r5810 := (r5809);
    r5811 := "0";
    null;
    r5812 := (r5811);
    r5813 := "0";
    null;
    r5814 := (r5813);
    r5815 := "0";
    null;
    r5816 := (r5815);
    r5817 := "1";
    null;
    r5818 := (r5817);
    r5819 := "0";
    null;
    r5820 := (r5819);
    r5821 := "1";
    null;
    r5822 := (r5821);
    r5823 := "1";
    null;
    r5824 := (r5823);
    r5825 := "0";
    null;
    r5826 := (r5825);
    r5827 := "1";
    null;
    r5828 := (r5827);
    r5829 := "1";
    null;
    r5830 := (r5829);
    r5831 := "1";
    null;
    r5832 := (r5831);
    r5833 := "0";
    null;
    r5834 := (r5833);
    r5835 := "0";
    null;
    r5836 := (r5835);
    r5837 := "0";
    null;
    r5838 := (r5837);
    r5839 := "0";
    null;
    r5840 := (r5839);
    r5776 := (r5778 & r5780 & r5782 & r5784 & r5786 & r5788 & r5790 & r5792 & r5794 & r5796 & r5798 & r5800 & r5802 & r5804 & r5806 & r5808 & r5810 & r5812 & r5814 & r5816 & r5818 & r5820 & r5822 & r5824 & r5826 & r5828 & r5830 & r5832 & r5834 & r5836 & r5838 & r5840);
    return r5776;
  end rewire_MetaprogrammingRWwc24b8b70_5775;
  function rewire_MetaprogrammingRWwa81a664b_5706 return std_logic_vector
  is
    variable r5771 : std_logic_vector(0 to 0) := (others => '0');
    variable r5770 : std_logic_vector(0 to 0) := (others => '0');
    variable r5769 : std_logic_vector(0 to 0) := (others => '0');
    variable r5768 : std_logic_vector(0 to 0) := (others => '0');
    variable r5767 : std_logic_vector(0 to 0) := (others => '0');
    variable r5766 : std_logic_vector(0 to 0) := (others => '0');
    variable r5765 : std_logic_vector(0 to 0) := (others => '0');
    variable r5764 : std_logic_vector(0 to 0) := (others => '0');
    variable r5763 : std_logic_vector(0 to 0) := (others => '0');
    variable r5762 : std_logic_vector(0 to 0) := (others => '0');
    variable r5761 : std_logic_vector(0 to 0) := (others => '0');
    variable r5760 : std_logic_vector(0 to 0) := (others => '0');
    variable r5759 : std_logic_vector(0 to 0) := (others => '0');
    variable r5758 : std_logic_vector(0 to 0) := (others => '0');
    variable r5757 : std_logic_vector(0 to 0) := (others => '0');
    variable r5756 : std_logic_vector(0 to 0) := (others => '0');
    variable r5755 : std_logic_vector(0 to 0) := (others => '0');
    variable r5754 : std_logic_vector(0 to 0) := (others => '0');
    variable r5753 : std_logic_vector(0 to 0) := (others => '0');
    variable r5752 : std_logic_vector(0 to 0) := (others => '0');
    variable r5751 : std_logic_vector(0 to 0) := (others => '0');
    variable r5750 : std_logic_vector(0 to 0) := (others => '0');
    variable r5749 : std_logic_vector(0 to 0) := (others => '0');
    variable r5748 : std_logic_vector(0 to 0) := (others => '0');
    variable r5747 : std_logic_vector(0 to 0) := (others => '0');
    variable r5746 : std_logic_vector(0 to 0) := (others => '0');
    variable r5745 : std_logic_vector(0 to 0) := (others => '0');
    variable r5744 : std_logic_vector(0 to 0) := (others => '0');
    variable r5743 : std_logic_vector(0 to 0) := (others => '0');
    variable r5742 : std_logic_vector(0 to 0) := (others => '0');
    variable r5741 : std_logic_vector(0 to 0) := (others => '0');
    variable r5740 : std_logic_vector(0 to 0) := (others => '0');
    variable r5739 : std_logic_vector(0 to 0) := (others => '0');
    variable r5738 : std_logic_vector(0 to 0) := (others => '0');
    variable r5737 : std_logic_vector(0 to 0) := (others => '0');
    variable r5736 : std_logic_vector(0 to 0) := (others => '0');
    variable r5735 : std_logic_vector(0 to 0) := (others => '0');
    variable r5734 : std_logic_vector(0 to 0) := (others => '0');
    variable r5733 : std_logic_vector(0 to 0) := (others => '0');
    variable r5732 : std_logic_vector(0 to 0) := (others => '0');
    variable r5731 : std_logic_vector(0 to 0) := (others => '0');
    variable r5730 : std_logic_vector(0 to 0) := (others => '0');
    variable r5729 : std_logic_vector(0 to 0) := (others => '0');
    variable r5728 : std_logic_vector(0 to 0) := (others => '0');
    variable r5727 : std_logic_vector(0 to 0) := (others => '0');
    variable r5726 : std_logic_vector(0 to 0) := (others => '0');
    variable r5725 : std_logic_vector(0 to 0) := (others => '0');
    variable r5724 : std_logic_vector(0 to 0) := (others => '0');
    variable r5723 : std_logic_vector(0 to 0) := (others => '0');
    variable r5722 : std_logic_vector(0 to 0) := (others => '0');
    variable r5721 : std_logic_vector(0 to 0) := (others => '0');
    variable r5720 : std_logic_vector(0 to 0) := (others => '0');
    variable r5719 : std_logic_vector(0 to 0) := (others => '0');
    variable r5718 : std_logic_vector(0 to 0) := (others => '0');
    variable r5717 : std_logic_vector(0 to 0) := (others => '0');
    variable r5716 : std_logic_vector(0 to 0) := (others => '0');
    variable r5715 : std_logic_vector(0 to 0) := (others => '0');
    variable r5714 : std_logic_vector(0 to 0) := (others => '0');
    variable r5713 : std_logic_vector(0 to 0) := (others => '0');
    variable r5712 : std_logic_vector(0 to 0) := (others => '0');
    variable r5711 : std_logic_vector(0 to 0) := (others => '0');
    variable r5710 : std_logic_vector(0 to 0) := (others => '0');
    variable r5709 : std_logic_vector(0 to 0) := (others => '0');
    variable r5708 : std_logic_vector(0 to 0) := (others => '0');
    variable r5707 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r5708 := "1";
    null;
    r5709 := (r5708);
    r5710 := "0";
    null;
    r5711 := (r5710);
    r5712 := "1";
    null;
    r5713 := (r5712);
    r5714 := "0";
    null;
    r5715 := (r5714);
    r5716 := "1";
    null;
    r5717 := (r5716);
    r5718 := "0";
    null;
    r5719 := (r5718);
    r5720 := "0";
    null;
    r5721 := (r5720);
    r5722 := "0";
    null;
    r5723 := (r5722);
    r5724 := "0";
    null;
    r5725 := (r5724);
    r5726 := "0";
    null;
    r5727 := (r5726);
    r5728 := "0";
    null;
    r5729 := (r5728);
    r5730 := "1";
    null;
    r5731 := (r5730);
    r5732 := "1";
    null;
    r5733 := (r5732);
    r5734 := "0";
    null;
    r5735 := (r5734);
    r5736 := "1";
    null;
    r5737 := (r5736);
    r5738 := "0";
    null;
    r5739 := (r5738);
    r5740 := "0";
    null;
    r5741 := (r5740);
    r5742 := "1";
    null;
    r5743 := (r5742);
    r5744 := "1";
    null;
    r5745 := (r5744);
    r5746 := "0";
    null;
    r5747 := (r5746);
    r5748 := "0";
    null;
    r5749 := (r5748);
    r5750 := "1";
    null;
    r5751 := (r5750);
    r5752 := "1";
    null;
    r5753 := (r5752);
    r5754 := "0";
    null;
    r5755 := (r5754);
    r5756 := "0";
    null;
    r5757 := (r5756);
    r5758 := "1";
    null;
    r5759 := (r5758);
    r5760 := "0";
    null;
    r5761 := (r5760);
    r5762 := "0";
    null;
    r5763 := (r5762);
    r5764 := "1";
    null;
    r5765 := (r5764);
    r5766 := "0";
    null;
    r5767 := (r5766);
    r5768 := "1";
    null;
    r5769 := (r5768);
    r5770 := "1";
    null;
    r5771 := (r5770);
    r5707 := (r5709 & r5711 & r5713 & r5715 & r5717 & r5719 & r5721 & r5723 & r5725 & r5727 & r5729 & r5731 & r5733 & r5735 & r5737 & r5739 & r5741 & r5743 & r5745 & r5747 & r5749 & r5751 & r5753 & r5755 & r5757 & r5759 & r5761 & r5763 & r5765 & r5767 & r5769 & r5771);
    return r5707;
  end rewire_MetaprogrammingRWwa81a664b_5706;
  function rewire_MetaprogrammingRWwa2bfe8a1_5637 return std_logic_vector
  is
    variable r5702 : std_logic_vector(0 to 0) := (others => '0');
    variable r5701 : std_logic_vector(0 to 0) := (others => '0');
    variable r5700 : std_logic_vector(0 to 0) := (others => '0');
    variable r5699 : std_logic_vector(0 to 0) := (others => '0');
    variable r5698 : std_logic_vector(0 to 0) := (others => '0');
    variable r5697 : std_logic_vector(0 to 0) := (others => '0');
    variable r5696 : std_logic_vector(0 to 0) := (others => '0');
    variable r5695 : std_logic_vector(0 to 0) := (others => '0');
    variable r5694 : std_logic_vector(0 to 0) := (others => '0');
    variable r5693 : std_logic_vector(0 to 0) := (others => '0');
    variable r5692 : std_logic_vector(0 to 0) := (others => '0');
    variable r5691 : std_logic_vector(0 to 0) := (others => '0');
    variable r5690 : std_logic_vector(0 to 0) := (others => '0');
    variable r5689 : std_logic_vector(0 to 0) := (others => '0');
    variable r5688 : std_logic_vector(0 to 0) := (others => '0');
    variable r5687 : std_logic_vector(0 to 0) := (others => '0');
    variable r5686 : std_logic_vector(0 to 0) := (others => '0');
    variable r5685 : std_logic_vector(0 to 0) := (others => '0');
    variable r5684 : std_logic_vector(0 to 0) := (others => '0');
    variable r5683 : std_logic_vector(0 to 0) := (others => '0');
    variable r5682 : std_logic_vector(0 to 0) := (others => '0');
    variable r5681 : std_logic_vector(0 to 0) := (others => '0');
    variable r5680 : std_logic_vector(0 to 0) := (others => '0');
    variable r5679 : std_logic_vector(0 to 0) := (others => '0');
    variable r5678 : std_logic_vector(0 to 0) := (others => '0');
    variable r5677 : std_logic_vector(0 to 0) := (others => '0');
    variable r5676 : std_logic_vector(0 to 0) := (others => '0');
    variable r5675 : std_logic_vector(0 to 0) := (others => '0');
    variable r5674 : std_logic_vector(0 to 0) := (others => '0');
    variable r5673 : std_logic_vector(0 to 0) := (others => '0');
    variable r5672 : std_logic_vector(0 to 0) := (others => '0');
    variable r5671 : std_logic_vector(0 to 0) := (others => '0');
    variable r5670 : std_logic_vector(0 to 0) := (others => '0');
    variable r5669 : std_logic_vector(0 to 0) := (others => '0');
    variable r5668 : std_logic_vector(0 to 0) := (others => '0');
    variable r5667 : std_logic_vector(0 to 0) := (others => '0');
    variable r5666 : std_logic_vector(0 to 0) := (others => '0');
    variable r5665 : std_logic_vector(0 to 0) := (others => '0');
    variable r5664 : std_logic_vector(0 to 0) := (others => '0');
    variable r5663 : std_logic_vector(0 to 0) := (others => '0');
    variable r5662 : std_logic_vector(0 to 0) := (others => '0');
    variable r5661 : std_logic_vector(0 to 0) := (others => '0');
    variable r5660 : std_logic_vector(0 to 0) := (others => '0');
    variable r5659 : std_logic_vector(0 to 0) := (others => '0');
    variable r5658 : std_logic_vector(0 to 0) := (others => '0');
    variable r5657 : std_logic_vector(0 to 0) := (others => '0');
    variable r5656 : std_logic_vector(0 to 0) := (others => '0');
    variable r5655 : std_logic_vector(0 to 0) := (others => '0');
    variable r5654 : std_logic_vector(0 to 0) := (others => '0');
    variable r5653 : std_logic_vector(0 to 0) := (others => '0');
    variable r5652 : std_logic_vector(0 to 0) := (others => '0');
    variable r5651 : std_logic_vector(0 to 0) := (others => '0');
    variable r5650 : std_logic_vector(0 to 0) := (others => '0');
    variable r5649 : std_logic_vector(0 to 0) := (others => '0');
    variable r5648 : std_logic_vector(0 to 0) := (others => '0');
    variable r5647 : std_logic_vector(0 to 0) := (others => '0');
    variable r5646 : std_logic_vector(0 to 0) := (others => '0');
    variable r5645 : std_logic_vector(0 to 0) := (others => '0');
    variable r5644 : std_logic_vector(0 to 0) := (others => '0');
    variable r5643 : std_logic_vector(0 to 0) := (others => '0');
    variable r5642 : std_logic_vector(0 to 0) := (others => '0');
    variable r5641 : std_logic_vector(0 to 0) := (others => '0');
    variable r5640 : std_logic_vector(0 to 0) := (others => '0');
    variable r5639 : std_logic_vector(0 to 0) := (others => '0');
    variable r5638 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r5639 := "1";
    null;
    r5640 := (r5639);
    r5641 := "0";
    null;
    r5642 := (r5641);
    r5643 := "1";
    null;
    r5644 := (r5643);
    r5645 := "0";
    null;
    r5646 := (r5645);
    r5647 := "0";
    null;
    r5648 := (r5647);
    r5649 := "0";
    null;
    r5650 := (r5649);
    r5651 := "1";
    null;
    r5652 := (r5651);
    r5653 := "0";
    null;
    r5654 := (r5653);
    r5655 := "1";
    null;
    r5656 := (r5655);
    r5657 := "0";
    null;
    r5658 := (r5657);
    r5659 := "1";
    null;
    r5660 := (r5659);
    r5661 := "1";
    null;
    r5662 := (r5661);
    r5663 := "1";
    null;
    r5664 := (r5663);
    r5665 := "1";
    null;
    r5666 := (r5665);
    r5667 := "1";
    null;
    r5668 := (r5667);
    r5669 := "1";
    null;
    r5670 := (r5669);
    r5671 := "1";
    null;
    r5672 := (r5671);
    r5673 := "1";
    null;
    r5674 := (r5673);
    r5675 := "1";
    null;
    r5676 := (r5675);
    r5677 := "0";
    null;
    r5678 := (r5677);
    r5679 := "1";
    null;
    r5680 := (r5679);
    r5681 := "0";
    null;
    r5682 := (r5681);
    r5683 := "0";
    null;
    r5684 := (r5683);
    r5685 := "0";
    null;
    r5686 := (r5685);
    r5687 := "1";
    null;
    r5688 := (r5687);
    r5689 := "0";
    null;
    r5690 := (r5689);
    r5691 := "1";
    null;
    r5692 := (r5691);
    r5693 := "0";
    null;
    r5694 := (r5693);
    r5695 := "0";
    null;
    r5696 := (r5695);
    r5697 := "0";
    null;
    r5698 := (r5697);
    r5699 := "0";
    null;
    r5700 := (r5699);
    r5701 := "1";
    null;
    r5702 := (r5701);
    r5638 := (r5640 & r5642 & r5644 & r5646 & r5648 & r5650 & r5652 & r5654 & r5656 & r5658 & r5660 & r5662 & r5664 & r5666 & r5668 & r5670 & r5672 & r5674 & r5676 & r5678 & r5680 & r5682 & r5684 & r5686 & r5688 & r5690 & r5692 & r5694 & r5696 & r5698 & r5700 & r5702);
    return r5638;
  end rewire_MetaprogrammingRWwa2bfe8a1_5637;
  function rewire_MetaprogrammingRWw92722c85_5568 return std_logic_vector
  is
    variable r5633 : std_logic_vector(0 to 0) := (others => '0');
    variable r5632 : std_logic_vector(0 to 0) := (others => '0');
    variable r5631 : std_logic_vector(0 to 0) := (others => '0');
    variable r5630 : std_logic_vector(0 to 0) := (others => '0');
    variable r5629 : std_logic_vector(0 to 0) := (others => '0');
    variable r5628 : std_logic_vector(0 to 0) := (others => '0');
    variable r5627 : std_logic_vector(0 to 0) := (others => '0');
    variable r5626 : std_logic_vector(0 to 0) := (others => '0');
    variable r5625 : std_logic_vector(0 to 0) := (others => '0');
    variable r5624 : std_logic_vector(0 to 0) := (others => '0');
    variable r5623 : std_logic_vector(0 to 0) := (others => '0');
    variable r5622 : std_logic_vector(0 to 0) := (others => '0');
    variable r5621 : std_logic_vector(0 to 0) := (others => '0');
    variable r5620 : std_logic_vector(0 to 0) := (others => '0');
    variable r5619 : std_logic_vector(0 to 0) := (others => '0');
    variable r5618 : std_logic_vector(0 to 0) := (others => '0');
    variable r5617 : std_logic_vector(0 to 0) := (others => '0');
    variable r5616 : std_logic_vector(0 to 0) := (others => '0');
    variable r5615 : std_logic_vector(0 to 0) := (others => '0');
    variable r5614 : std_logic_vector(0 to 0) := (others => '0');
    variable r5613 : std_logic_vector(0 to 0) := (others => '0');
    variable r5612 : std_logic_vector(0 to 0) := (others => '0');
    variable r5611 : std_logic_vector(0 to 0) := (others => '0');
    variable r5610 : std_logic_vector(0 to 0) := (others => '0');
    variable r5609 : std_logic_vector(0 to 0) := (others => '0');
    variable r5608 : std_logic_vector(0 to 0) := (others => '0');
    variable r5607 : std_logic_vector(0 to 0) := (others => '0');
    variable r5606 : std_logic_vector(0 to 0) := (others => '0');
    variable r5605 : std_logic_vector(0 to 0) := (others => '0');
    variable r5604 : std_logic_vector(0 to 0) := (others => '0');
    variable r5603 : std_logic_vector(0 to 0) := (others => '0');
    variable r5602 : std_logic_vector(0 to 0) := (others => '0');
    variable r5601 : std_logic_vector(0 to 0) := (others => '0');
    variable r5600 : std_logic_vector(0 to 0) := (others => '0');
    variable r5599 : std_logic_vector(0 to 0) := (others => '0');
    variable r5598 : std_logic_vector(0 to 0) := (others => '0');
    variable r5597 : std_logic_vector(0 to 0) := (others => '0');
    variable r5596 : std_logic_vector(0 to 0) := (others => '0');
    variable r5595 : std_logic_vector(0 to 0) := (others => '0');
    variable r5594 : std_logic_vector(0 to 0) := (others => '0');
    variable r5593 : std_logic_vector(0 to 0) := (others => '0');
    variable r5592 : std_logic_vector(0 to 0) := (others => '0');
    variable r5591 : std_logic_vector(0 to 0) := (others => '0');
    variable r5590 : std_logic_vector(0 to 0) := (others => '0');
    variable r5589 : std_logic_vector(0 to 0) := (others => '0');
    variable r5588 : std_logic_vector(0 to 0) := (others => '0');
    variable r5587 : std_logic_vector(0 to 0) := (others => '0');
    variable r5586 : std_logic_vector(0 to 0) := (others => '0');
    variable r5585 : std_logic_vector(0 to 0) := (others => '0');
    variable r5584 : std_logic_vector(0 to 0) := (others => '0');
    variable r5583 : std_logic_vector(0 to 0) := (others => '0');
    variable r5582 : std_logic_vector(0 to 0) := (others => '0');
    variable r5581 : std_logic_vector(0 to 0) := (others => '0');
    variable r5580 : std_logic_vector(0 to 0) := (others => '0');
    variable r5579 : std_logic_vector(0 to 0) := (others => '0');
    variable r5578 : std_logic_vector(0 to 0) := (others => '0');
    variable r5577 : std_logic_vector(0 to 0) := (others => '0');
    variable r5576 : std_logic_vector(0 to 0) := (others => '0');
    variable r5575 : std_logic_vector(0 to 0) := (others => '0');
    variable r5574 : std_logic_vector(0 to 0) := (others => '0');
    variable r5573 : std_logic_vector(0 to 0) := (others => '0');
    variable r5572 : std_logic_vector(0 to 0) := (others => '0');
    variable r5571 : std_logic_vector(0 to 0) := (others => '0');
    variable r5570 : std_logic_vector(0 to 0) := (others => '0');
    variable r5569 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r5570 := "1";
    null;
    r5571 := (r5570);
    r5572 := "0";
    null;
    r5573 := (r5572);
    r5574 := "0";
    null;
    r5575 := (r5574);
    r5576 := "1";
    null;
    r5577 := (r5576);
    r5578 := "0";
    null;
    r5579 := (r5578);
    r5580 := "0";
    null;
    r5581 := (r5580);
    r5582 := "1";
    null;
    r5583 := (r5582);
    r5584 := "0";
    null;
    r5585 := (r5584);
    r5586 := "0";
    null;
    r5587 := (r5586);
    r5588 := "1";
    null;
    r5589 := (r5588);
    r5590 := "1";
    null;
    r5591 := (r5590);
    r5592 := "1";
    null;
    r5593 := (r5592);
    r5594 := "0";
    null;
    r5595 := (r5594);
    r5596 := "0";
    null;
    r5597 := (r5596);
    r5598 := "1";
    null;
    r5599 := (r5598);
    r5600 := "0";
    null;
    r5601 := (r5600);
    r5602 := "0";
    null;
    r5603 := (r5602);
    r5604 := "0";
    null;
    r5605 := (r5604);
    r5606 := "1";
    null;
    r5607 := (r5606);
    r5608 := "0";
    null;
    r5609 := (r5608);
    r5610 := "1";
    null;
    r5611 := (r5610);
    r5612 := "1";
    null;
    r5613 := (r5612);
    r5614 := "0";
    null;
    r5615 := (r5614);
    r5616 := "0";
    null;
    r5617 := (r5616);
    r5618 := "1";
    null;
    r5619 := (r5618);
    r5620 := "0";
    null;
    r5621 := (r5620);
    r5622 := "0";
    null;
    r5623 := (r5622);
    r5624 := "0";
    null;
    r5625 := (r5624);
    r5626 := "0";
    null;
    r5627 := (r5626);
    r5628 := "1";
    null;
    r5629 := (r5628);
    r5630 := "0";
    null;
    r5631 := (r5630);
    r5632 := "1";
    null;
    r5633 := (r5632);
    r5569 := (r5571 & r5573 & r5575 & r5577 & r5579 & r5581 & r5583 & r5585 & r5587 & r5589 & r5591 & r5593 & r5595 & r5597 & r5599 & r5601 & r5603 & r5605 & r5607 & r5609 & r5611 & r5613 & r5615 & r5617 & r5619 & r5621 & r5623 & r5625 & r5627 & r5629 & r5631 & r5633);
    return r5569;
  end rewire_MetaprogrammingRWw92722c85_5568;
  function rewire_MetaprogrammingRWw81c2c92e_5499 return std_logic_vector
  is
    variable r5564 : std_logic_vector(0 to 0) := (others => '0');
    variable r5563 : std_logic_vector(0 to 0) := (others => '0');
    variable r5562 : std_logic_vector(0 to 0) := (others => '0');
    variable r5561 : std_logic_vector(0 to 0) := (others => '0');
    variable r5560 : std_logic_vector(0 to 0) := (others => '0');
    variable r5559 : std_logic_vector(0 to 0) := (others => '0');
    variable r5558 : std_logic_vector(0 to 0) := (others => '0');
    variable r5557 : std_logic_vector(0 to 0) := (others => '0');
    variable r5556 : std_logic_vector(0 to 0) := (others => '0');
    variable r5555 : std_logic_vector(0 to 0) := (others => '0');
    variable r5554 : std_logic_vector(0 to 0) := (others => '0');
    variable r5553 : std_logic_vector(0 to 0) := (others => '0');
    variable r5552 : std_logic_vector(0 to 0) := (others => '0');
    variable r5551 : std_logic_vector(0 to 0) := (others => '0');
    variable r5550 : std_logic_vector(0 to 0) := (others => '0');
    variable r5549 : std_logic_vector(0 to 0) := (others => '0');
    variable r5548 : std_logic_vector(0 to 0) := (others => '0');
    variable r5547 : std_logic_vector(0 to 0) := (others => '0');
    variable r5546 : std_logic_vector(0 to 0) := (others => '0');
    variable r5545 : std_logic_vector(0 to 0) := (others => '0');
    variable r5544 : std_logic_vector(0 to 0) := (others => '0');
    variable r5543 : std_logic_vector(0 to 0) := (others => '0');
    variable r5542 : std_logic_vector(0 to 0) := (others => '0');
    variable r5541 : std_logic_vector(0 to 0) := (others => '0');
    variable r5540 : std_logic_vector(0 to 0) := (others => '0');
    variable r5539 : std_logic_vector(0 to 0) := (others => '0');
    variable r5538 : std_logic_vector(0 to 0) := (others => '0');
    variable r5537 : std_logic_vector(0 to 0) := (others => '0');
    variable r5536 : std_logic_vector(0 to 0) := (others => '0');
    variable r5535 : std_logic_vector(0 to 0) := (others => '0');
    variable r5534 : std_logic_vector(0 to 0) := (others => '0');
    variable r5533 : std_logic_vector(0 to 0) := (others => '0');
    variable r5532 : std_logic_vector(0 to 0) := (others => '0');
    variable r5531 : std_logic_vector(0 to 0) := (others => '0');
    variable r5530 : std_logic_vector(0 to 0) := (others => '0');
    variable r5529 : std_logic_vector(0 to 0) := (others => '0');
    variable r5528 : std_logic_vector(0 to 0) := (others => '0');
    variable r5527 : std_logic_vector(0 to 0) := (others => '0');
    variable r5526 : std_logic_vector(0 to 0) := (others => '0');
    variable r5525 : std_logic_vector(0 to 0) := (others => '0');
    variable r5524 : std_logic_vector(0 to 0) := (others => '0');
    variable r5523 : std_logic_vector(0 to 0) := (others => '0');
    variable r5522 : std_logic_vector(0 to 0) := (others => '0');
    variable r5521 : std_logic_vector(0 to 0) := (others => '0');
    variable r5520 : std_logic_vector(0 to 0) := (others => '0');
    variable r5519 : std_logic_vector(0 to 0) := (others => '0');
    variable r5518 : std_logic_vector(0 to 0) := (others => '0');
    variable r5517 : std_logic_vector(0 to 0) := (others => '0');
    variable r5516 : std_logic_vector(0 to 0) := (others => '0');
    variable r5515 : std_logic_vector(0 to 0) := (others => '0');
    variable r5514 : std_logic_vector(0 to 0) := (others => '0');
    variable r5513 : std_logic_vector(0 to 0) := (others => '0');
    variable r5512 : std_logic_vector(0 to 0) := (others => '0');
    variable r5511 : std_logic_vector(0 to 0) := (others => '0');
    variable r5510 : std_logic_vector(0 to 0) := (others => '0');
    variable r5509 : std_logic_vector(0 to 0) := (others => '0');
    variable r5508 : std_logic_vector(0 to 0) := (others => '0');
    variable r5507 : std_logic_vector(0 to 0) := (others => '0');
    variable r5506 : std_logic_vector(0 to 0) := (others => '0');
    variable r5505 : std_logic_vector(0 to 0) := (others => '0');
    variable r5504 : std_logic_vector(0 to 0) := (others => '0');
    variable r5503 : std_logic_vector(0 to 0) := (others => '0');
    variable r5502 : std_logic_vector(0 to 0) := (others => '0');
    variable r5501 : std_logic_vector(0 to 0) := (others => '0');
    variable r5500 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r5501 := "1";
    null;
    r5502 := (r5501);
    r5503 := "0";
    null;
    r5504 := (r5503);
    r5505 := "0";
    null;
    r5506 := (r5505);
    r5507 := "0";
    null;
    r5508 := (r5507);
    r5509 := "0";
    null;
    r5510 := (r5509);
    r5511 := "0";
    null;
    r5512 := (r5511);
    r5513 := "0";
    null;
    r5514 := (r5513);
    r5515 := "1";
    null;
    r5516 := (r5515);
    r5517 := "1";
    null;
    r5518 := (r5517);
    r5519 := "1";
    null;
    r5520 := (r5519);
    r5521 := "0";
    null;
    r5522 := (r5521);
    r5523 := "0";
    null;
    r5524 := (r5523);
    r5525 := "0";
    null;
    r5526 := (r5525);
    r5527 := "0";
    null;
    r5528 := (r5527);
    r5529 := "1";
    null;
    r5530 := (r5529);
    r5531 := "0";
    null;
    r5532 := (r5531);
    r5533 := "1";
    null;
    r5534 := (r5533);
    r5535 := "1";
    null;
    r5536 := (r5535);
    r5537 := "0";
    null;
    r5538 := (r5537);
    r5539 := "0";
    null;
    r5540 := (r5539);
    r5541 := "1";
    null;
    r5542 := (r5541);
    r5543 := "0";
    null;
    r5544 := (r5543);
    r5545 := "0";
    null;
    r5546 := (r5545);
    r5547 := "1";
    null;
    r5548 := (r5547);
    r5549 := "0";
    null;
    r5550 := (r5549);
    r5551 := "0";
    null;
    r5552 := (r5551);
    r5553 := "1";
    null;
    r5554 := (r5553);
    r5555 := "0";
    null;
    r5556 := (r5555);
    r5557 := "1";
    null;
    r5558 := (r5557);
    r5559 := "1";
    null;
    r5560 := (r5559);
    r5561 := "1";
    null;
    r5562 := (r5561);
    r5563 := "0";
    null;
    r5564 := (r5563);
    r5500 := (r5502 & r5504 & r5506 & r5508 & r5510 & r5512 & r5514 & r5516 & r5518 & r5520 & r5522 & r5524 & r5526 & r5528 & r5530 & r5532 & r5534 & r5536 & r5538 & r5540 & r5542 & r5544 & r5546 & r5548 & r5550 & r5552 & r5554 & r5556 & r5558 & r5560 & r5562 & r5564);
    return r5500;
  end rewire_MetaprogrammingRWw81c2c92e_5499;
  function rewire_MetaprogrammingRWw766a0abb_5430 return std_logic_vector
  is
    variable r5495 : std_logic_vector(0 to 0) := (others => '0');
    variable r5494 : std_logic_vector(0 to 0) := (others => '0');
    variable r5493 : std_logic_vector(0 to 0) := (others => '0');
    variable r5492 : std_logic_vector(0 to 0) := (others => '0');
    variable r5491 : std_logic_vector(0 to 0) := (others => '0');
    variable r5490 : std_logic_vector(0 to 0) := (others => '0');
    variable r5489 : std_logic_vector(0 to 0) := (others => '0');
    variable r5488 : std_logic_vector(0 to 0) := (others => '0');
    variable r5487 : std_logic_vector(0 to 0) := (others => '0');
    variable r5486 : std_logic_vector(0 to 0) := (others => '0');
    variable r5485 : std_logic_vector(0 to 0) := (others => '0');
    variable r5484 : std_logic_vector(0 to 0) := (others => '0');
    variable r5483 : std_logic_vector(0 to 0) := (others => '0');
    variable r5482 : std_logic_vector(0 to 0) := (others => '0');
    variable r5481 : std_logic_vector(0 to 0) := (others => '0');
    variable r5480 : std_logic_vector(0 to 0) := (others => '0');
    variable r5479 : std_logic_vector(0 to 0) := (others => '0');
    variable r5478 : std_logic_vector(0 to 0) := (others => '0');
    variable r5477 : std_logic_vector(0 to 0) := (others => '0');
    variable r5476 : std_logic_vector(0 to 0) := (others => '0');
    variable r5475 : std_logic_vector(0 to 0) := (others => '0');
    variable r5474 : std_logic_vector(0 to 0) := (others => '0');
    variable r5473 : std_logic_vector(0 to 0) := (others => '0');
    variable r5472 : std_logic_vector(0 to 0) := (others => '0');
    variable r5471 : std_logic_vector(0 to 0) := (others => '0');
    variable r5470 : std_logic_vector(0 to 0) := (others => '0');
    variable r5469 : std_logic_vector(0 to 0) := (others => '0');
    variable r5468 : std_logic_vector(0 to 0) := (others => '0');
    variable r5467 : std_logic_vector(0 to 0) := (others => '0');
    variable r5466 : std_logic_vector(0 to 0) := (others => '0');
    variable r5465 : std_logic_vector(0 to 0) := (others => '0');
    variable r5464 : std_logic_vector(0 to 0) := (others => '0');
    variable r5463 : std_logic_vector(0 to 0) := (others => '0');
    variable r5462 : std_logic_vector(0 to 0) := (others => '0');
    variable r5461 : std_logic_vector(0 to 0) := (others => '0');
    variable r5460 : std_logic_vector(0 to 0) := (others => '0');
    variable r5459 : std_logic_vector(0 to 0) := (others => '0');
    variable r5458 : std_logic_vector(0 to 0) := (others => '0');
    variable r5457 : std_logic_vector(0 to 0) := (others => '0');
    variable r5456 : std_logic_vector(0 to 0) := (others => '0');
    variable r5455 : std_logic_vector(0 to 0) := (others => '0');
    variable r5454 : std_logic_vector(0 to 0) := (others => '0');
    variable r5453 : std_logic_vector(0 to 0) := (others => '0');
    variable r5452 : std_logic_vector(0 to 0) := (others => '0');
    variable r5451 : std_logic_vector(0 to 0) := (others => '0');
    variable r5450 : std_logic_vector(0 to 0) := (others => '0');
    variable r5449 : std_logic_vector(0 to 0) := (others => '0');
    variable r5448 : std_logic_vector(0 to 0) := (others => '0');
    variable r5447 : std_logic_vector(0 to 0) := (others => '0');
    variable r5446 : std_logic_vector(0 to 0) := (others => '0');
    variable r5445 : std_logic_vector(0 to 0) := (others => '0');
    variable r5444 : std_logic_vector(0 to 0) := (others => '0');
    variable r5443 : std_logic_vector(0 to 0) := (others => '0');
    variable r5442 : std_logic_vector(0 to 0) := (others => '0');
    variable r5441 : std_logic_vector(0 to 0) := (others => '0');
    variable r5440 : std_logic_vector(0 to 0) := (others => '0');
    variable r5439 : std_logic_vector(0 to 0) := (others => '0');
    variable r5438 : std_logic_vector(0 to 0) := (others => '0');
    variable r5437 : std_logic_vector(0 to 0) := (others => '0');
    variable r5436 : std_logic_vector(0 to 0) := (others => '0');
    variable r5435 : std_logic_vector(0 to 0) := (others => '0');
    variable r5434 : std_logic_vector(0 to 0) := (others => '0');
    variable r5433 : std_logic_vector(0 to 0) := (others => '0');
    variable r5432 : std_logic_vector(0 to 0) := (others => '0');
    variable r5431 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r5432 := "0";
    null;
    r5433 := (r5432);
    r5434 := "1";
    null;
    r5435 := (r5434);
    r5436 := "1";
    null;
    r5437 := (r5436);
    r5438 := "1";
    null;
    r5439 := (r5438);
    r5440 := "0";
    null;
    r5441 := (r5440);
    r5442 := "1";
    null;
    r5443 := (r5442);
    r5444 := "1";
    null;
    r5445 := (r5444);
    r5446 := "0";
    null;
    r5447 := (r5446);
    r5448 := "0";
    null;
    r5449 := (r5448);
    r5450 := "1";
    null;
    r5451 := (r5450);
    r5452 := "1";
    null;
    r5453 := (r5452);
    r5454 := "0";
    null;
    r5455 := (r5454);
    r5456 := "1";
    null;
    r5457 := (r5456);
    r5458 := "0";
    null;
    r5459 := (r5458);
    r5460 := "1";
    null;
    r5461 := (r5460);
    r5462 := "0";
    null;
    r5463 := (r5462);
    r5464 := "0";
    null;
    r5465 := (r5464);
    r5466 := "0";
    null;
    r5467 := (r5466);
    r5468 := "0";
    null;
    r5469 := (r5468);
    r5470 := "0";
    null;
    r5471 := (r5470);
    r5472 := "1";
    null;
    r5473 := (r5472);
    r5474 := "0";
    null;
    r5475 := (r5474);
    r5476 := "1";
    null;
    r5477 := (r5476);
    r5478 := "0";
    null;
    r5479 := (r5478);
    r5480 := "1";
    null;
    r5481 := (r5480);
    r5482 := "0";
    null;
    r5483 := (r5482);
    r5484 := "1";
    null;
    r5485 := (r5484);
    r5486 := "1";
    null;
    r5487 := (r5486);
    r5488 := "1";
    null;
    r5489 := (r5488);
    r5490 := "0";
    null;
    r5491 := (r5490);
    r5492 := "1";
    null;
    r5493 := (r5492);
    r5494 := "1";
    null;
    r5495 := (r5494);
    r5431 := (r5433 & r5435 & r5437 & r5439 & r5441 & r5443 & r5445 & r5447 & r5449 & r5451 & r5453 & r5455 & r5457 & r5459 & r5461 & r5463 & r5465 & r5467 & r5469 & r5471 & r5473 & r5475 & r5477 & r5479 & r5481 & r5483 & r5485 & r5487 & r5489 & r5491 & r5493 & r5495);
    return r5431;
  end rewire_MetaprogrammingRWw766a0abb_5430;
  function rewire_MetaprogrammingRWw650a7354_5361 return std_logic_vector
  is
    variable r5426 : std_logic_vector(0 to 0) := (others => '0');
    variable r5425 : std_logic_vector(0 to 0) := (others => '0');
    variable r5424 : std_logic_vector(0 to 0) := (others => '0');
    variable r5423 : std_logic_vector(0 to 0) := (others => '0');
    variable r5422 : std_logic_vector(0 to 0) := (others => '0');
    variable r5421 : std_logic_vector(0 to 0) := (others => '0');
    variable r5420 : std_logic_vector(0 to 0) := (others => '0');
    variable r5419 : std_logic_vector(0 to 0) := (others => '0');
    variable r5418 : std_logic_vector(0 to 0) := (others => '0');
    variable r5417 : std_logic_vector(0 to 0) := (others => '0');
    variable r5416 : std_logic_vector(0 to 0) := (others => '0');
    variable r5415 : std_logic_vector(0 to 0) := (others => '0');
    variable r5414 : std_logic_vector(0 to 0) := (others => '0');
    variable r5413 : std_logic_vector(0 to 0) := (others => '0');
    variable r5412 : std_logic_vector(0 to 0) := (others => '0');
    variable r5411 : std_logic_vector(0 to 0) := (others => '0');
    variable r5410 : std_logic_vector(0 to 0) := (others => '0');
    variable r5409 : std_logic_vector(0 to 0) := (others => '0');
    variable r5408 : std_logic_vector(0 to 0) := (others => '0');
    variable r5407 : std_logic_vector(0 to 0) := (others => '0');
    variable r5406 : std_logic_vector(0 to 0) := (others => '0');
    variable r5405 : std_logic_vector(0 to 0) := (others => '0');
    variable r5404 : std_logic_vector(0 to 0) := (others => '0');
    variable r5403 : std_logic_vector(0 to 0) := (others => '0');
    variable r5402 : std_logic_vector(0 to 0) := (others => '0');
    variable r5401 : std_logic_vector(0 to 0) := (others => '0');
    variable r5400 : std_logic_vector(0 to 0) := (others => '0');
    variable r5399 : std_logic_vector(0 to 0) := (others => '0');
    variable r5398 : std_logic_vector(0 to 0) := (others => '0');
    variable r5397 : std_logic_vector(0 to 0) := (others => '0');
    variable r5396 : std_logic_vector(0 to 0) := (others => '0');
    variable r5395 : std_logic_vector(0 to 0) := (others => '0');
    variable r5394 : std_logic_vector(0 to 0) := (others => '0');
    variable r5393 : std_logic_vector(0 to 0) := (others => '0');
    variable r5392 : std_logic_vector(0 to 0) := (others => '0');
    variable r5391 : std_logic_vector(0 to 0) := (others => '0');
    variable r5390 : std_logic_vector(0 to 0) := (others => '0');
    variable r5389 : std_logic_vector(0 to 0) := (others => '0');
    variable r5388 : std_logic_vector(0 to 0) := (others => '0');
    variable r5387 : std_logic_vector(0 to 0) := (others => '0');
    variable r5386 : std_logic_vector(0 to 0) := (others => '0');
    variable r5385 : std_logic_vector(0 to 0) := (others => '0');
    variable r5384 : std_logic_vector(0 to 0) := (others => '0');
    variable r5383 : std_logic_vector(0 to 0) := (others => '0');
    variable r5382 : std_logic_vector(0 to 0) := (others => '0');
    variable r5381 : std_logic_vector(0 to 0) := (others => '0');
    variable r5380 : std_logic_vector(0 to 0) := (others => '0');
    variable r5379 : std_logic_vector(0 to 0) := (others => '0');
    variable r5378 : std_logic_vector(0 to 0) := (others => '0');
    variable r5377 : std_logic_vector(0 to 0) := (others => '0');
    variable r5376 : std_logic_vector(0 to 0) := (others => '0');
    variable r5375 : std_logic_vector(0 to 0) := (others => '0');
    variable r5374 : std_logic_vector(0 to 0) := (others => '0');
    variable r5373 : std_logic_vector(0 to 0) := (others => '0');
    variable r5372 : std_logic_vector(0 to 0) := (others => '0');
    variable r5371 : std_logic_vector(0 to 0) := (others => '0');
    variable r5370 : std_logic_vector(0 to 0) := (others => '0');
    variable r5369 : std_logic_vector(0 to 0) := (others => '0');
    variable r5368 : std_logic_vector(0 to 0) := (others => '0');
    variable r5367 : std_logic_vector(0 to 0) := (others => '0');
    variable r5366 : std_logic_vector(0 to 0) := (others => '0');
    variable r5365 : std_logic_vector(0 to 0) := (others => '0');
    variable r5364 : std_logic_vector(0 to 0) := (others => '0');
    variable r5363 : std_logic_vector(0 to 0) := (others => '0');
    variable r5362 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r5363 := "0";
    null;
    r5364 := (r5363);
    r5365 := "1";
    null;
    r5366 := (r5365);
    r5367 := "1";
    null;
    r5368 := (r5367);
    r5369 := "0";
    null;
    r5370 := (r5369);
    r5371 := "0";
    null;
    r5372 := (r5371);
    r5373 := "1";
    null;
    r5374 := (r5373);
    r5375 := "0";
    null;
    r5376 := (r5375);
    r5377 := "1";
    null;
    r5378 := (r5377);
    r5379 := "0";
    null;
    r5380 := (r5379);
    r5381 := "0";
    null;
    r5382 := (r5381);
    r5383 := "0";
    null;
    r5384 := (r5383);
    r5385 := "0";
    null;
    r5386 := (r5385);
    r5387 := "1";
    null;
    r5388 := (r5387);
    r5389 := "0";
    null;
    r5390 := (r5389);
    r5391 := "1";
    null;
    r5392 := (r5391);
    r5393 := "0";
    null;
    r5394 := (r5393);
    r5395 := "0";
    null;
    r5396 := (r5395);
    r5397 := "1";
    null;
    r5398 := (r5397);
    r5399 := "1";
    null;
    r5400 := (r5399);
    r5401 := "1";
    null;
    r5402 := (r5401);
    r5403 := "0";
    null;
    r5404 := (r5403);
    r5405 := "0";
    null;
    r5406 := (r5405);
    r5407 := "1";
    null;
    r5408 := (r5407);
    r5409 := "1";
    null;
    r5410 := (r5409);
    r5411 := "0";
    null;
    r5412 := (r5411);
    r5413 := "1";
    null;
    r5414 := (r5413);
    r5415 := "0";
    null;
    r5416 := (r5415);
    r5417 := "1";
    null;
    r5418 := (r5417);
    r5419 := "0";
    null;
    r5420 := (r5419);
    r5421 := "1";
    null;
    r5422 := (r5421);
    r5423 := "0";
    null;
    r5424 := (r5423);
    r5425 := "0";
    null;
    r5426 := (r5425);
    r5362 := (r5364 & r5366 & r5368 & r5370 & r5372 & r5374 & r5376 & r5378 & r5380 & r5382 & r5384 & r5386 & r5388 & r5390 & r5392 & r5394 & r5396 & r5398 & r5400 & r5402 & r5404 & r5406 & r5408 & r5410 & r5412 & r5414 & r5416 & r5418 & r5420 & r5422 & r5424 & r5426);
    return r5362;
  end rewire_MetaprogrammingRWw650a7354_5361;
  function rewire_MetaprogrammingRWw53380d13_5292 return std_logic_vector
  is
    variable r5357 : std_logic_vector(0 to 0) := (others => '0');
    variable r5356 : std_logic_vector(0 to 0) := (others => '0');
    variable r5355 : std_logic_vector(0 to 0) := (others => '0');
    variable r5354 : std_logic_vector(0 to 0) := (others => '0');
    variable r5353 : std_logic_vector(0 to 0) := (others => '0');
    variable r5352 : std_logic_vector(0 to 0) := (others => '0');
    variable r5351 : std_logic_vector(0 to 0) := (others => '0');
    variable r5350 : std_logic_vector(0 to 0) := (others => '0');
    variable r5349 : std_logic_vector(0 to 0) := (others => '0');
    variable r5348 : std_logic_vector(0 to 0) := (others => '0');
    variable r5347 : std_logic_vector(0 to 0) := (others => '0');
    variable r5346 : std_logic_vector(0 to 0) := (others => '0');
    variable r5345 : std_logic_vector(0 to 0) := (others => '0');
    variable r5344 : std_logic_vector(0 to 0) := (others => '0');
    variable r5343 : std_logic_vector(0 to 0) := (others => '0');
    variable r5342 : std_logic_vector(0 to 0) := (others => '0');
    variable r5341 : std_logic_vector(0 to 0) := (others => '0');
    variable r5340 : std_logic_vector(0 to 0) := (others => '0');
    variable r5339 : std_logic_vector(0 to 0) := (others => '0');
    variable r5338 : std_logic_vector(0 to 0) := (others => '0');
    variable r5337 : std_logic_vector(0 to 0) := (others => '0');
    variable r5336 : std_logic_vector(0 to 0) := (others => '0');
    variable r5335 : std_logic_vector(0 to 0) := (others => '0');
    variable r5334 : std_logic_vector(0 to 0) := (others => '0');
    variable r5333 : std_logic_vector(0 to 0) := (others => '0');
    variable r5332 : std_logic_vector(0 to 0) := (others => '0');
    variable r5331 : std_logic_vector(0 to 0) := (others => '0');
    variable r5330 : std_logic_vector(0 to 0) := (others => '0');
    variable r5329 : std_logic_vector(0 to 0) := (others => '0');
    variable r5328 : std_logic_vector(0 to 0) := (others => '0');
    variable r5327 : std_logic_vector(0 to 0) := (others => '0');
    variable r5326 : std_logic_vector(0 to 0) := (others => '0');
    variable r5325 : std_logic_vector(0 to 0) := (others => '0');
    variable r5324 : std_logic_vector(0 to 0) := (others => '0');
    variable r5323 : std_logic_vector(0 to 0) := (others => '0');
    variable r5322 : std_logic_vector(0 to 0) := (others => '0');
    variable r5321 : std_logic_vector(0 to 0) := (others => '0');
    variable r5320 : std_logic_vector(0 to 0) := (others => '0');
    variable r5319 : std_logic_vector(0 to 0) := (others => '0');
    variable r5318 : std_logic_vector(0 to 0) := (others => '0');
    variable r5317 : std_logic_vector(0 to 0) := (others => '0');
    variable r5316 : std_logic_vector(0 to 0) := (others => '0');
    variable r5315 : std_logic_vector(0 to 0) := (others => '0');
    variable r5314 : std_logic_vector(0 to 0) := (others => '0');
    variable r5313 : std_logic_vector(0 to 0) := (others => '0');
    variable r5312 : std_logic_vector(0 to 0) := (others => '0');
    variable r5311 : std_logic_vector(0 to 0) := (others => '0');
    variable r5310 : std_logic_vector(0 to 0) := (others => '0');
    variable r5309 : std_logic_vector(0 to 0) := (others => '0');
    variable r5308 : std_logic_vector(0 to 0) := (others => '0');
    variable r5307 : std_logic_vector(0 to 0) := (others => '0');
    variable r5306 : std_logic_vector(0 to 0) := (others => '0');
    variable r5305 : std_logic_vector(0 to 0) := (others => '0');
    variable r5304 : std_logic_vector(0 to 0) := (others => '0');
    variable r5303 : std_logic_vector(0 to 0) := (others => '0');
    variable r5302 : std_logic_vector(0 to 0) := (others => '0');
    variable r5301 : std_logic_vector(0 to 0) := (others => '0');
    variable r5300 : std_logic_vector(0 to 0) := (others => '0');
    variable r5299 : std_logic_vector(0 to 0) := (others => '0');
    variable r5298 : std_logic_vector(0 to 0) := (others => '0');
    variable r5297 : std_logic_vector(0 to 0) := (others => '0');
    variable r5296 : std_logic_vector(0 to 0) := (others => '0');
    variable r5295 : std_logic_vector(0 to 0) := (others => '0');
    variable r5294 : std_logic_vector(0 to 0) := (others => '0');
    variable r5293 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r5294 := "0";
    null;
    r5295 := (r5294);
    r5296 := "1";
    null;
    r5297 := (r5296);
    r5298 := "0";
    null;
    r5299 := (r5298);
    r5300 := "1";
    null;
    r5301 := (r5300);
    r5302 := "0";
    null;
    r5303 := (r5302);
    r5304 := "0";
    null;
    r5305 := (r5304);
    r5306 := "1";
    null;
    r5307 := (r5306);
    r5308 := "1";
    null;
    r5309 := (r5308);
    r5310 := "0";
    null;
    r5311 := (r5310);
    r5312 := "0";
    null;
    r5313 := (r5312);
    r5314 := "1";
    null;
    r5315 := (r5314);
    r5316 := "1";
    null;
    r5317 := (r5316);
    r5318 := "1";
    null;
    r5319 := (r5318);
    r5320 := "0";
    null;
    r5321 := (r5320);
    r5322 := "0";
    null;
    r5323 := (r5322);
    r5324 := "0";
    null;
    r5325 := (r5324);
    r5326 := "0";
    null;
    r5327 := (r5326);
    r5328 := "0";
    null;
    r5329 := (r5328);
    r5330 := "0";
    null;
    r5331 := (r5330);
    r5332 := "0";
    null;
    r5333 := (r5332);
    r5334 := "1";
    null;
    r5335 := (r5334);
    r5336 := "1";
    null;
    r5337 := (r5336);
    r5338 := "0";
    null;
    r5339 := (r5338);
    r5340 := "1";
    null;
    r5341 := (r5340);
    r5342 := "0";
    null;
    r5343 := (r5342);
    r5344 := "0";
    null;
    r5345 := (r5344);
    r5346 := "0";
    null;
    r5347 := (r5346);
    r5348 := "1";
    null;
    r5349 := (r5348);
    r5350 := "0";
    null;
    r5351 := (r5350);
    r5352 := "0";
    null;
    r5353 := (r5352);
    r5354 := "1";
    null;
    r5355 := (r5354);
    r5356 := "1";
    null;
    r5357 := (r5356);
    r5293 := (r5295 & r5297 & r5299 & r5301 & r5303 & r5305 & r5307 & r5309 & r5311 & r5313 & r5315 & r5317 & r5319 & r5321 & r5323 & r5325 & r5327 & r5329 & r5331 & r5333 & r5335 & r5337 & r5339 & r5341 & r5343 & r5345 & r5347 & r5349 & r5351 & r5353 & r5355 & r5357);
    return r5293;
  end rewire_MetaprogrammingRWw53380d13_5292;
  function rewire_MetaprogrammingRWw4d2c6dfc_5223 return std_logic_vector
  is
    variable r5288 : std_logic_vector(0 to 0) := (others => '0');
    variable r5287 : std_logic_vector(0 to 0) := (others => '0');
    variable r5286 : std_logic_vector(0 to 0) := (others => '0');
    variable r5285 : std_logic_vector(0 to 0) := (others => '0');
    variable r5284 : std_logic_vector(0 to 0) := (others => '0');
    variable r5283 : std_logic_vector(0 to 0) := (others => '0');
    variable r5282 : std_logic_vector(0 to 0) := (others => '0');
    variable r5281 : std_logic_vector(0 to 0) := (others => '0');
    variable r5280 : std_logic_vector(0 to 0) := (others => '0');
    variable r5279 : std_logic_vector(0 to 0) := (others => '0');
    variable r5278 : std_logic_vector(0 to 0) := (others => '0');
    variable r5277 : std_logic_vector(0 to 0) := (others => '0');
    variable r5276 : std_logic_vector(0 to 0) := (others => '0');
    variable r5275 : std_logic_vector(0 to 0) := (others => '0');
    variable r5274 : std_logic_vector(0 to 0) := (others => '0');
    variable r5273 : std_logic_vector(0 to 0) := (others => '0');
    variable r5272 : std_logic_vector(0 to 0) := (others => '0');
    variable r5271 : std_logic_vector(0 to 0) := (others => '0');
    variable r5270 : std_logic_vector(0 to 0) := (others => '0');
    variable r5269 : std_logic_vector(0 to 0) := (others => '0');
    variable r5268 : std_logic_vector(0 to 0) := (others => '0');
    variable r5267 : std_logic_vector(0 to 0) := (others => '0');
    variable r5266 : std_logic_vector(0 to 0) := (others => '0');
    variable r5265 : std_logic_vector(0 to 0) := (others => '0');
    variable r5264 : std_logic_vector(0 to 0) := (others => '0');
    variable r5263 : std_logic_vector(0 to 0) := (others => '0');
    variable r5262 : std_logic_vector(0 to 0) := (others => '0');
    variable r5261 : std_logic_vector(0 to 0) := (others => '0');
    variable r5260 : std_logic_vector(0 to 0) := (others => '0');
    variable r5259 : std_logic_vector(0 to 0) := (others => '0');
    variable r5258 : std_logic_vector(0 to 0) := (others => '0');
    variable r5257 : std_logic_vector(0 to 0) := (others => '0');
    variable r5256 : std_logic_vector(0 to 0) := (others => '0');
    variable r5255 : std_logic_vector(0 to 0) := (others => '0');
    variable r5254 : std_logic_vector(0 to 0) := (others => '0');
    variable r5253 : std_logic_vector(0 to 0) := (others => '0');
    variable r5252 : std_logic_vector(0 to 0) := (others => '0');
    variable r5251 : std_logic_vector(0 to 0) := (others => '0');
    variable r5250 : std_logic_vector(0 to 0) := (others => '0');
    variable r5249 : std_logic_vector(0 to 0) := (others => '0');
    variable r5248 : std_logic_vector(0 to 0) := (others => '0');
    variable r5247 : std_logic_vector(0 to 0) := (others => '0');
    variable r5246 : std_logic_vector(0 to 0) := (others => '0');
    variable r5245 : std_logic_vector(0 to 0) := (others => '0');
    variable r5244 : std_logic_vector(0 to 0) := (others => '0');
    variable r5243 : std_logic_vector(0 to 0) := (others => '0');
    variable r5242 : std_logic_vector(0 to 0) := (others => '0');
    variable r5241 : std_logic_vector(0 to 0) := (others => '0');
    variable r5240 : std_logic_vector(0 to 0) := (others => '0');
    variable r5239 : std_logic_vector(0 to 0) := (others => '0');
    variable r5238 : std_logic_vector(0 to 0) := (others => '0');
    variable r5237 : std_logic_vector(0 to 0) := (others => '0');
    variable r5236 : std_logic_vector(0 to 0) := (others => '0');
    variable r5235 : std_logic_vector(0 to 0) := (others => '0');
    variable r5234 : std_logic_vector(0 to 0) := (others => '0');
    variable r5233 : std_logic_vector(0 to 0) := (others => '0');
    variable r5232 : std_logic_vector(0 to 0) := (others => '0');
    variable r5231 : std_logic_vector(0 to 0) := (others => '0');
    variable r5230 : std_logic_vector(0 to 0) := (others => '0');
    variable r5229 : std_logic_vector(0 to 0) := (others => '0');
    variable r5228 : std_logic_vector(0 to 0) := (others => '0');
    variable r5227 : std_logic_vector(0 to 0) := (others => '0');
    variable r5226 : std_logic_vector(0 to 0) := (others => '0');
    variable r5225 : std_logic_vector(0 to 0) := (others => '0');
    variable r5224 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r5225 := "0";
    null;
    r5226 := (r5225);
    r5227 := "1";
    null;
    r5228 := (r5227);
    r5229 := "0";
    null;
    r5230 := (r5229);
    r5231 := "0";
    null;
    r5232 := (r5231);
    r5233 := "1";
    null;
    r5234 := (r5233);
    r5235 := "1";
    null;
    r5236 := (r5235);
    r5237 := "0";
    null;
    r5238 := (r5237);
    r5239 := "1";
    null;
    r5240 := (r5239);
    r5241 := "0";
    null;
    r5242 := (r5241);
    r5243 := "0";
    null;
    r5244 := (r5243);
    r5245 := "1";
    null;
    r5246 := (r5245);
    r5247 := "0";
    null;
    r5248 := (r5247);
    r5249 := "1";
    null;
    r5250 := (r5249);
    r5251 := "1";
    null;
    r5252 := (r5251);
    r5253 := "0";
    null;
    r5254 := (r5253);
    r5255 := "0";
    null;
    r5256 := (r5255);
    r5257 := "0";
    null;
    r5258 := (r5257);
    r5259 := "1";
    null;
    r5260 := (r5259);
    r5261 := "1";
    null;
    r5262 := (r5261);
    r5263 := "0";
    null;
    r5264 := (r5263);
    r5265 := "1";
    null;
    r5266 := (r5265);
    r5267 := "1";
    null;
    r5268 := (r5267);
    r5269 := "0";
    null;
    r5270 := (r5269);
    r5271 := "1";
    null;
    r5272 := (r5271);
    r5273 := "1";
    null;
    r5274 := (r5273);
    r5275 := "1";
    null;
    r5276 := (r5275);
    r5277 := "1";
    null;
    r5278 := (r5277);
    r5279 := "1";
    null;
    r5280 := (r5279);
    r5281 := "1";
    null;
    r5282 := (r5281);
    r5283 := "1";
    null;
    r5284 := (r5283);
    r5285 := "0";
    null;
    r5286 := (r5285);
    r5287 := "0";
    null;
    r5288 := (r5287);
    r5224 := (r5226 & r5228 & r5230 & r5232 & r5234 & r5236 & r5238 & r5240 & r5242 & r5244 & r5246 & r5248 & r5250 & r5252 & r5254 & r5256 & r5258 & r5260 & r5262 & r5264 & r5266 & r5268 & r5270 & r5272 & r5274 & r5276 & r5278 & r5280 & r5282 & r5284 & r5286 & r5288);
    return r5224;
  end rewire_MetaprogrammingRWw4d2c6dfc_5223;
  function rewire_MetaprogrammingRWw2e1b2138_5154 return std_logic_vector
  is
    variable r5219 : std_logic_vector(0 to 0) := (others => '0');
    variable r5218 : std_logic_vector(0 to 0) := (others => '0');
    variable r5217 : std_logic_vector(0 to 0) := (others => '0');
    variable r5216 : std_logic_vector(0 to 0) := (others => '0');
    variable r5215 : std_logic_vector(0 to 0) := (others => '0');
    variable r5214 : std_logic_vector(0 to 0) := (others => '0');
    variable r5213 : std_logic_vector(0 to 0) := (others => '0');
    variable r5212 : std_logic_vector(0 to 0) := (others => '0');
    variable r5211 : std_logic_vector(0 to 0) := (others => '0');
    variable r5210 : std_logic_vector(0 to 0) := (others => '0');
    variable r5209 : std_logic_vector(0 to 0) := (others => '0');
    variable r5208 : std_logic_vector(0 to 0) := (others => '0');
    variable r5207 : std_logic_vector(0 to 0) := (others => '0');
    variable r5206 : std_logic_vector(0 to 0) := (others => '0');
    variable r5205 : std_logic_vector(0 to 0) := (others => '0');
    variable r5204 : std_logic_vector(0 to 0) := (others => '0');
    variable r5203 : std_logic_vector(0 to 0) := (others => '0');
    variable r5202 : std_logic_vector(0 to 0) := (others => '0');
    variable r5201 : std_logic_vector(0 to 0) := (others => '0');
    variable r5200 : std_logic_vector(0 to 0) := (others => '0');
    variable r5199 : std_logic_vector(0 to 0) := (others => '0');
    variable r5198 : std_logic_vector(0 to 0) := (others => '0');
    variable r5197 : std_logic_vector(0 to 0) := (others => '0');
    variable r5196 : std_logic_vector(0 to 0) := (others => '0');
    variable r5195 : std_logic_vector(0 to 0) := (others => '0');
    variable r5194 : std_logic_vector(0 to 0) := (others => '0');
    variable r5193 : std_logic_vector(0 to 0) := (others => '0');
    variable r5192 : std_logic_vector(0 to 0) := (others => '0');
    variable r5191 : std_logic_vector(0 to 0) := (others => '0');
    variable r5190 : std_logic_vector(0 to 0) := (others => '0');
    variable r5189 : std_logic_vector(0 to 0) := (others => '0');
    variable r5188 : std_logic_vector(0 to 0) := (others => '0');
    variable r5187 : std_logic_vector(0 to 0) := (others => '0');
    variable r5186 : std_logic_vector(0 to 0) := (others => '0');
    variable r5185 : std_logic_vector(0 to 0) := (others => '0');
    variable r5184 : std_logic_vector(0 to 0) := (others => '0');
    variable r5183 : std_logic_vector(0 to 0) := (others => '0');
    variable r5182 : std_logic_vector(0 to 0) := (others => '0');
    variable r5181 : std_logic_vector(0 to 0) := (others => '0');
    variable r5180 : std_logic_vector(0 to 0) := (others => '0');
    variable r5179 : std_logic_vector(0 to 0) := (others => '0');
    variable r5178 : std_logic_vector(0 to 0) := (others => '0');
    variable r5177 : std_logic_vector(0 to 0) := (others => '0');
    variable r5176 : std_logic_vector(0 to 0) := (others => '0');
    variable r5175 : std_logic_vector(0 to 0) := (others => '0');
    variable r5174 : std_logic_vector(0 to 0) := (others => '0');
    variable r5173 : std_logic_vector(0 to 0) := (others => '0');
    variable r5172 : std_logic_vector(0 to 0) := (others => '0');
    variable r5171 : std_logic_vector(0 to 0) := (others => '0');
    variable r5170 : std_logic_vector(0 to 0) := (others => '0');
    variable r5169 : std_logic_vector(0 to 0) := (others => '0');
    variable r5168 : std_logic_vector(0 to 0) := (others => '0');
    variable r5167 : std_logic_vector(0 to 0) := (others => '0');
    variable r5166 : std_logic_vector(0 to 0) := (others => '0');
    variable r5165 : std_logic_vector(0 to 0) := (others => '0');
    variable r5164 : std_logic_vector(0 to 0) := (others => '0');
    variable r5163 : std_logic_vector(0 to 0) := (others => '0');
    variable r5162 : std_logic_vector(0 to 0) := (others => '0');
    variable r5161 : std_logic_vector(0 to 0) := (others => '0');
    variable r5160 : std_logic_vector(0 to 0) := (others => '0');
    variable r5159 : std_logic_vector(0 to 0) := (others => '0');
    variable r5158 : std_logic_vector(0 to 0) := (others => '0');
    variable r5157 : std_logic_vector(0 to 0) := (others => '0');
    variable r5156 : std_logic_vector(0 to 0) := (others => '0');
    variable r5155 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r5156 := "0";
    null;
    r5157 := (r5156);
    r5158 := "0";
    null;
    r5159 := (r5158);
    r5160 := "1";
    null;
    r5161 := (r5160);
    r5162 := "0";
    null;
    r5163 := (r5162);
    r5164 := "1";
    null;
    r5165 := (r5164);
    r5166 := "1";
    null;
    r5167 := (r5166);
    r5168 := "1";
    null;
    r5169 := (r5168);
    r5170 := "0";
    null;
    r5171 := (r5170);
    r5172 := "0";
    null;
    r5173 := (r5172);
    r5174 := "0";
    null;
    r5175 := (r5174);
    r5176 := "0";
    null;
    r5177 := (r5176);
    r5178 := "1";
    null;
    r5179 := (r5178);
    r5180 := "1";
    null;
    r5181 := (r5180);
    r5182 := "0";
    null;
    r5183 := (r5182);
    r5184 := "1";
    null;
    r5185 := (r5184);
    r5186 := "1";
    null;
    r5187 := (r5186);
    r5188 := "0";
    null;
    r5189 := (r5188);
    r5190 := "0";
    null;
    r5191 := (r5190);
    r5192 := "1";
    null;
    r5193 := (r5192);
    r5194 := "0";
    null;
    r5195 := (r5194);
    r5196 := "0";
    null;
    r5197 := (r5196);
    r5198 := "0";
    null;
    r5199 := (r5198);
    r5200 := "0";
    null;
    r5201 := (r5200);
    r5202 := "1";
    null;
    r5203 := (r5202);
    r5204 := "0";
    null;
    r5205 := (r5204);
    r5206 := "0";
    null;
    r5207 := (r5206);
    r5208 := "1";
    null;
    r5209 := (r5208);
    r5210 := "1";
    null;
    r5211 := (r5210);
    r5212 := "1";
    null;
    r5213 := (r5212);
    r5214 := "0";
    null;
    r5215 := (r5214);
    r5216 := "0";
    null;
    r5217 := (r5216);
    r5218 := "0";
    null;
    r5219 := (r5218);
    r5155 := (r5157 & r5159 & r5161 & r5163 & r5165 & r5167 & r5169 & r5171 & r5173 & r5175 & r5177 & r5179 & r5181 & r5183 & r5185 & r5187 & r5189 & r5191 & r5193 & r5195 & r5197 & r5199 & r5201 & r5203 & r5205 & r5207 & r5209 & r5211 & r5213 & r5215 & r5217 & r5219);
    return r5155;
  end rewire_MetaprogrammingRWw2e1b2138_5154;
  function rewire_MetaprogrammingRWw27b70a85_5085 return std_logic_vector
  is
    variable r5150 : std_logic_vector(0 to 0) := (others => '0');
    variable r5149 : std_logic_vector(0 to 0) := (others => '0');
    variable r5148 : std_logic_vector(0 to 0) := (others => '0');
    variable r5147 : std_logic_vector(0 to 0) := (others => '0');
    variable r5146 : std_logic_vector(0 to 0) := (others => '0');
    variable r5145 : std_logic_vector(0 to 0) := (others => '0');
    variable r5144 : std_logic_vector(0 to 0) := (others => '0');
    variable r5143 : std_logic_vector(0 to 0) := (others => '0');
    variable r5142 : std_logic_vector(0 to 0) := (others => '0');
    variable r5141 : std_logic_vector(0 to 0) := (others => '0');
    variable r5140 : std_logic_vector(0 to 0) := (others => '0');
    variable r5139 : std_logic_vector(0 to 0) := (others => '0');
    variable r5138 : std_logic_vector(0 to 0) := (others => '0');
    variable r5137 : std_logic_vector(0 to 0) := (others => '0');
    variable r5136 : std_logic_vector(0 to 0) := (others => '0');
    variable r5135 : std_logic_vector(0 to 0) := (others => '0');
    variable r5134 : std_logic_vector(0 to 0) := (others => '0');
    variable r5133 : std_logic_vector(0 to 0) := (others => '0');
    variable r5132 : std_logic_vector(0 to 0) := (others => '0');
    variable r5131 : std_logic_vector(0 to 0) := (others => '0');
    variable r5130 : std_logic_vector(0 to 0) := (others => '0');
    variable r5129 : std_logic_vector(0 to 0) := (others => '0');
    variable r5128 : std_logic_vector(0 to 0) := (others => '0');
    variable r5127 : std_logic_vector(0 to 0) := (others => '0');
    variable r5126 : std_logic_vector(0 to 0) := (others => '0');
    variable r5125 : std_logic_vector(0 to 0) := (others => '0');
    variable r5124 : std_logic_vector(0 to 0) := (others => '0');
    variable r5123 : std_logic_vector(0 to 0) := (others => '0');
    variable r5122 : std_logic_vector(0 to 0) := (others => '0');
    variable r5121 : std_logic_vector(0 to 0) := (others => '0');
    variable r5120 : std_logic_vector(0 to 0) := (others => '0');
    variable r5119 : std_logic_vector(0 to 0) := (others => '0');
    variable r5118 : std_logic_vector(0 to 0) := (others => '0');
    variable r5117 : std_logic_vector(0 to 0) := (others => '0');
    variable r5116 : std_logic_vector(0 to 0) := (others => '0');
    variable r5115 : std_logic_vector(0 to 0) := (others => '0');
    variable r5114 : std_logic_vector(0 to 0) := (others => '0');
    variable r5113 : std_logic_vector(0 to 0) := (others => '0');
    variable r5112 : std_logic_vector(0 to 0) := (others => '0');
    variable r5111 : std_logic_vector(0 to 0) := (others => '0');
    variable r5110 : std_logic_vector(0 to 0) := (others => '0');
    variable r5109 : std_logic_vector(0 to 0) := (others => '0');
    variable r5108 : std_logic_vector(0 to 0) := (others => '0');
    variable r5107 : std_logic_vector(0 to 0) := (others => '0');
    variable r5106 : std_logic_vector(0 to 0) := (others => '0');
    variable r5105 : std_logic_vector(0 to 0) := (others => '0');
    variable r5104 : std_logic_vector(0 to 0) := (others => '0');
    variable r5103 : std_logic_vector(0 to 0) := (others => '0');
    variable r5102 : std_logic_vector(0 to 0) := (others => '0');
    variable r5101 : std_logic_vector(0 to 0) := (others => '0');
    variable r5100 : std_logic_vector(0 to 0) := (others => '0');
    variable r5099 : std_logic_vector(0 to 0) := (others => '0');
    variable r5098 : std_logic_vector(0 to 0) := (others => '0');
    variable r5097 : std_logic_vector(0 to 0) := (others => '0');
    variable r5096 : std_logic_vector(0 to 0) := (others => '0');
    variable r5095 : std_logic_vector(0 to 0) := (others => '0');
    variable r5094 : std_logic_vector(0 to 0) := (others => '0');
    variable r5093 : std_logic_vector(0 to 0) := (others => '0');
    variable r5092 : std_logic_vector(0 to 0) := (others => '0');
    variable r5091 : std_logic_vector(0 to 0) := (others => '0');
    variable r5090 : std_logic_vector(0 to 0) := (others => '0');
    variable r5089 : std_logic_vector(0 to 0) := (others => '0');
    variable r5088 : std_logic_vector(0 to 0) := (others => '0');
    variable r5087 : std_logic_vector(0 to 0) := (others => '0');
    variable r5086 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r5087 := "0";
    null;
    r5088 := (r5087);
    r5089 := "0";
    null;
    r5090 := (r5089);
    r5091 := "1";
    null;
    r5092 := (r5091);
    r5093 := "0";
    null;
    r5094 := (r5093);
    r5095 := "0";
    null;
    r5096 := (r5095);
    r5097 := "1";
    null;
    r5098 := (r5097);
    r5099 := "1";
    null;
    r5100 := (r5099);
    r5101 := "1";
    null;
    r5102 := (r5101);
    r5103 := "1";
    null;
    r5104 := (r5103);
    r5105 := "0";
    null;
    r5106 := (r5105);
    r5107 := "1";
    null;
    r5108 := (r5107);
    r5109 := "1";
    null;
    r5110 := (r5109);
    r5111 := "0";
    null;
    r5112 := (r5111);
    r5113 := "1";
    null;
    r5114 := (r5113);
    r5115 := "1";
    null;
    r5116 := (r5115);
    r5117 := "1";
    null;
    r5118 := (r5117);
    r5119 := "0";
    null;
    r5120 := (r5119);
    r5121 := "0";
    null;
    r5122 := (r5121);
    r5123 := "0";
    null;
    r5124 := (r5123);
    r5125 := "0";
    null;
    r5126 := (r5125);
    r5127 := "1";
    null;
    r5128 := (r5127);
    r5129 := "0";
    null;
    r5130 := (r5129);
    r5131 := "1";
    null;
    r5132 := (r5131);
    r5133 := "0";
    null;
    r5134 := (r5133);
    r5135 := "1";
    null;
    r5136 := (r5135);
    r5137 := "0";
    null;
    r5138 := (r5137);
    r5139 := "0";
    null;
    r5140 := (r5139);
    r5141 := "0";
    null;
    r5142 := (r5141);
    r5143 := "0";
    null;
    r5144 := (r5143);
    r5145 := "1";
    null;
    r5146 := (r5145);
    r5147 := "0";
    null;
    r5148 := (r5147);
    r5149 := "1";
    null;
    r5150 := (r5149);
    r5086 := (r5088 & r5090 & r5092 & r5094 & r5096 & r5098 & r5100 & r5102 & r5104 & r5106 & r5108 & r5110 & r5112 & r5114 & r5116 & r5118 & r5120 & r5122 & r5124 & r5126 & r5128 & r5130 & r5132 & r5134 & r5136 & r5138 & r5140 & r5142 & r5144 & r5146 & r5148 & r5150);
    return r5086;
  end rewire_MetaprogrammingRWw27b70a85_5085;
  function rewire_MetaprogrammingRWw14292967_5016 return std_logic_vector
  is
    variable r5081 : std_logic_vector(0 to 0) := (others => '0');
    variable r5080 : std_logic_vector(0 to 0) := (others => '0');
    variable r5079 : std_logic_vector(0 to 0) := (others => '0');
    variable r5078 : std_logic_vector(0 to 0) := (others => '0');
    variable r5077 : std_logic_vector(0 to 0) := (others => '0');
    variable r5076 : std_logic_vector(0 to 0) := (others => '0');
    variable r5075 : std_logic_vector(0 to 0) := (others => '0');
    variable r5074 : std_logic_vector(0 to 0) := (others => '0');
    variable r5073 : std_logic_vector(0 to 0) := (others => '0');
    variable r5072 : std_logic_vector(0 to 0) := (others => '0');
    variable r5071 : std_logic_vector(0 to 0) := (others => '0');
    variable r5070 : std_logic_vector(0 to 0) := (others => '0');
    variable r5069 : std_logic_vector(0 to 0) := (others => '0');
    variable r5068 : std_logic_vector(0 to 0) := (others => '0');
    variable r5067 : std_logic_vector(0 to 0) := (others => '0');
    variable r5066 : std_logic_vector(0 to 0) := (others => '0');
    variable r5065 : std_logic_vector(0 to 0) := (others => '0');
    variable r5064 : std_logic_vector(0 to 0) := (others => '0');
    variable r5063 : std_logic_vector(0 to 0) := (others => '0');
    variable r5062 : std_logic_vector(0 to 0) := (others => '0');
    variable r5061 : std_logic_vector(0 to 0) := (others => '0');
    variable r5060 : std_logic_vector(0 to 0) := (others => '0');
    variable r5059 : std_logic_vector(0 to 0) := (others => '0');
    variable r5058 : std_logic_vector(0 to 0) := (others => '0');
    variable r5057 : std_logic_vector(0 to 0) := (others => '0');
    variable r5056 : std_logic_vector(0 to 0) := (others => '0');
    variable r5055 : std_logic_vector(0 to 0) := (others => '0');
    variable r5054 : std_logic_vector(0 to 0) := (others => '0');
    variable r5053 : std_logic_vector(0 to 0) := (others => '0');
    variable r5052 : std_logic_vector(0 to 0) := (others => '0');
    variable r5051 : std_logic_vector(0 to 0) := (others => '0');
    variable r5050 : std_logic_vector(0 to 0) := (others => '0');
    variable r5049 : std_logic_vector(0 to 0) := (others => '0');
    variable r5048 : std_logic_vector(0 to 0) := (others => '0');
    variable r5047 : std_logic_vector(0 to 0) := (others => '0');
    variable r5046 : std_logic_vector(0 to 0) := (others => '0');
    variable r5045 : std_logic_vector(0 to 0) := (others => '0');
    variable r5044 : std_logic_vector(0 to 0) := (others => '0');
    variable r5043 : std_logic_vector(0 to 0) := (others => '0');
    variable r5042 : std_logic_vector(0 to 0) := (others => '0');
    variable r5041 : std_logic_vector(0 to 0) := (others => '0');
    variable r5040 : std_logic_vector(0 to 0) := (others => '0');
    variable r5039 : std_logic_vector(0 to 0) := (others => '0');
    variable r5038 : std_logic_vector(0 to 0) := (others => '0');
    variable r5037 : std_logic_vector(0 to 0) := (others => '0');
    variable r5036 : std_logic_vector(0 to 0) := (others => '0');
    variable r5035 : std_logic_vector(0 to 0) := (others => '0');
    variable r5034 : std_logic_vector(0 to 0) := (others => '0');
    variable r5033 : std_logic_vector(0 to 0) := (others => '0');
    variable r5032 : std_logic_vector(0 to 0) := (others => '0');
    variable r5031 : std_logic_vector(0 to 0) := (others => '0');
    variable r5030 : std_logic_vector(0 to 0) := (others => '0');
    variable r5029 : std_logic_vector(0 to 0) := (others => '0');
    variable r5028 : std_logic_vector(0 to 0) := (others => '0');
    variable r5027 : std_logic_vector(0 to 0) := (others => '0');
    variable r5026 : std_logic_vector(0 to 0) := (others => '0');
    variable r5025 : std_logic_vector(0 to 0) := (others => '0');
    variable r5024 : std_logic_vector(0 to 0) := (others => '0');
    variable r5023 : std_logic_vector(0 to 0) := (others => '0');
    variable r5022 : std_logic_vector(0 to 0) := (others => '0');
    variable r5021 : std_logic_vector(0 to 0) := (others => '0');
    variable r5020 : std_logic_vector(0 to 0) := (others => '0');
    variable r5019 : std_logic_vector(0 to 0) := (others => '0');
    variable r5018 : std_logic_vector(0 to 0) := (others => '0');
    variable r5017 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r5018 := "0";
    null;
    r5019 := (r5018);
    r5020 := "0";
    null;
    r5021 := (r5020);
    r5022 := "0";
    null;
    r5023 := (r5022);
    r5024 := "1";
    null;
    r5025 := (r5024);
    r5026 := "0";
    null;
    r5027 := (r5026);
    r5028 := "1";
    null;
    r5029 := (r5028);
    r5030 := "0";
    null;
    r5031 := (r5030);
    r5032 := "0";
    null;
    r5033 := (r5032);
    r5034 := "0";
    null;
    r5035 := (r5034);
    r5036 := "0";
    null;
    r5037 := (r5036);
    r5038 := "1";
    null;
    r5039 := (r5038);
    r5040 := "0";
    null;
    r5041 := (r5040);
    r5042 := "1";
    null;
    r5043 := (r5042);
    r5044 := "0";
    null;
    r5045 := (r5044);
    r5046 := "0";
    null;
    r5047 := (r5046);
    r5048 := "1";
    null;
    r5049 := (r5048);
    r5050 := "0";
    null;
    r5051 := (r5050);
    r5052 := "0";
    null;
    r5053 := (r5052);
    r5054 := "1";
    null;
    r5055 := (r5054);
    r5056 := "0";
    null;
    r5057 := (r5056);
    r5058 := "1";
    null;
    r5059 := (r5058);
    r5060 := "0";
    null;
    r5061 := (r5060);
    r5062 := "0";
    null;
    r5063 := (r5062);
    r5064 := "1";
    null;
    r5065 := (r5064);
    r5066 := "0";
    null;
    r5067 := (r5066);
    r5068 := "1";
    null;
    r5069 := (r5068);
    r5070 := "1";
    null;
    r5071 := (r5070);
    r5072 := "0";
    null;
    r5073 := (r5072);
    r5074 := "0";
    null;
    r5075 := (r5074);
    r5076 := "1";
    null;
    r5077 := (r5076);
    r5078 := "1";
    null;
    r5079 := (r5078);
    r5080 := "1";
    null;
    r5081 := (r5080);
    r5017 := (r5019 & r5021 & r5023 & r5025 & r5027 & r5029 & r5031 & r5033 & r5035 & r5037 & r5039 & r5041 & r5043 & r5045 & r5047 & r5049 & r5051 & r5053 & r5055 & r5057 & r5059 & r5061 & r5063 & r5065 & r5067 & r5069 & r5071 & r5073 & r5075 & r5077 & r5079 & r5081);
    return r5017;
  end rewire_MetaprogrammingRWw14292967_5016;
  function rewire_MetaprogrammingRWw06ca6351_4947 return std_logic_vector
  is
    variable r5012 : std_logic_vector(0 to 0) := (others => '0');
    variable r5011 : std_logic_vector(0 to 0) := (others => '0');
    variable r5010 : std_logic_vector(0 to 0) := (others => '0');
    variable r5009 : std_logic_vector(0 to 0) := (others => '0');
    variable r5008 : std_logic_vector(0 to 0) := (others => '0');
    variable r5007 : std_logic_vector(0 to 0) := (others => '0');
    variable r5006 : std_logic_vector(0 to 0) := (others => '0');
    variable r5005 : std_logic_vector(0 to 0) := (others => '0');
    variable r5004 : std_logic_vector(0 to 0) := (others => '0');
    variable r5003 : std_logic_vector(0 to 0) := (others => '0');
    variable r5002 : std_logic_vector(0 to 0) := (others => '0');
    variable r5001 : std_logic_vector(0 to 0) := (others => '0');
    variable r5000 : std_logic_vector(0 to 0) := (others => '0');
    variable r4999 : std_logic_vector(0 to 0) := (others => '0');
    variable r4998 : std_logic_vector(0 to 0) := (others => '0');
    variable r4997 : std_logic_vector(0 to 0) := (others => '0');
    variable r4996 : std_logic_vector(0 to 0) := (others => '0');
    variable r4995 : std_logic_vector(0 to 0) := (others => '0');
    variable r4994 : std_logic_vector(0 to 0) := (others => '0');
    variable r4993 : std_logic_vector(0 to 0) := (others => '0');
    variable r4992 : std_logic_vector(0 to 0) := (others => '0');
    variable r4991 : std_logic_vector(0 to 0) := (others => '0');
    variable r4990 : std_logic_vector(0 to 0) := (others => '0');
    variable r4989 : std_logic_vector(0 to 0) := (others => '0');
    variable r4988 : std_logic_vector(0 to 0) := (others => '0');
    variable r4987 : std_logic_vector(0 to 0) := (others => '0');
    variable r4986 : std_logic_vector(0 to 0) := (others => '0');
    variable r4985 : std_logic_vector(0 to 0) := (others => '0');
    variable r4984 : std_logic_vector(0 to 0) := (others => '0');
    variable r4983 : std_logic_vector(0 to 0) := (others => '0');
    variable r4982 : std_logic_vector(0 to 0) := (others => '0');
    variable r4981 : std_logic_vector(0 to 0) := (others => '0');
    variable r4980 : std_logic_vector(0 to 0) := (others => '0');
    variable r4979 : std_logic_vector(0 to 0) := (others => '0');
    variable r4978 : std_logic_vector(0 to 0) := (others => '0');
    variable r4977 : std_logic_vector(0 to 0) := (others => '0');
    variable r4976 : std_logic_vector(0 to 0) := (others => '0');
    variable r4975 : std_logic_vector(0 to 0) := (others => '0');
    variable r4974 : std_logic_vector(0 to 0) := (others => '0');
    variable r4973 : std_logic_vector(0 to 0) := (others => '0');
    variable r4972 : std_logic_vector(0 to 0) := (others => '0');
    variable r4971 : std_logic_vector(0 to 0) := (others => '0');
    variable r4970 : std_logic_vector(0 to 0) := (others => '0');
    variable r4969 : std_logic_vector(0 to 0) := (others => '0');
    variable r4968 : std_logic_vector(0 to 0) := (others => '0');
    variable r4967 : std_logic_vector(0 to 0) := (others => '0');
    variable r4966 : std_logic_vector(0 to 0) := (others => '0');
    variable r4965 : std_logic_vector(0 to 0) := (others => '0');
    variable r4964 : std_logic_vector(0 to 0) := (others => '0');
    variable r4963 : std_logic_vector(0 to 0) := (others => '0');
    variable r4962 : std_logic_vector(0 to 0) := (others => '0');
    variable r4961 : std_logic_vector(0 to 0) := (others => '0');
    variable r4960 : std_logic_vector(0 to 0) := (others => '0');
    variable r4959 : std_logic_vector(0 to 0) := (others => '0');
    variable r4958 : std_logic_vector(0 to 0) := (others => '0');
    variable r4957 : std_logic_vector(0 to 0) := (others => '0');
    variable r4956 : std_logic_vector(0 to 0) := (others => '0');
    variable r4955 : std_logic_vector(0 to 0) := (others => '0');
    variable r4954 : std_logic_vector(0 to 0) := (others => '0');
    variable r4953 : std_logic_vector(0 to 0) := (others => '0');
    variable r4952 : std_logic_vector(0 to 0) := (others => '0');
    variable r4951 : std_logic_vector(0 to 0) := (others => '0');
    variable r4950 : std_logic_vector(0 to 0) := (others => '0');
    variable r4949 : std_logic_vector(0 to 0) := (others => '0');
    variable r4948 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r4949 := "0";
    null;
    r4950 := (r4949);
    r4951 := "0";
    null;
    r4952 := (r4951);
    r4953 := "0";
    null;
    r4954 := (r4953);
    r4955 := "0";
    null;
    r4956 := (r4955);
    r4957 := "0";
    null;
    r4958 := (r4957);
    r4959 := "1";
    null;
    r4960 := (r4959);
    r4961 := "1";
    null;
    r4962 := (r4961);
    r4963 := "0";
    null;
    r4964 := (r4963);
    r4965 := "1";
    null;
    r4966 := (r4965);
    r4967 := "1";
    null;
    r4968 := (r4967);
    r4969 := "0";
    null;
    r4970 := (r4969);
    r4971 := "0";
    null;
    r4972 := (r4971);
    r4973 := "1";
    null;
    r4974 := (r4973);
    r4975 := "0";
    null;
    r4976 := (r4975);
    r4977 := "1";
    null;
    r4978 := (r4977);
    r4979 := "0";
    null;
    r4980 := (r4979);
    r4981 := "0";
    null;
    r4982 := (r4981);
    r4983 := "1";
    null;
    r4984 := (r4983);
    r4985 := "1";
    null;
    r4986 := (r4985);
    r4987 := "0";
    null;
    r4988 := (r4987);
    r4989 := "0";
    null;
    r4990 := (r4989);
    r4991 := "0";
    null;
    r4992 := (r4991);
    r4993 := "1";
    null;
    r4994 := (r4993);
    r4995 := "1";
    null;
    r4996 := (r4995);
    r4997 := "0";
    null;
    r4998 := (r4997);
    r4999 := "1";
    null;
    r5000 := (r4999);
    r5001 := "0";
    null;
    r5002 := (r5001);
    r5003 := "1";
    null;
    r5004 := (r5003);
    r5005 := "0";
    null;
    r5006 := (r5005);
    r5007 := "0";
    null;
    r5008 := (r5007);
    r5009 := "0";
    null;
    r5010 := (r5009);
    r5011 := "1";
    null;
    r5012 := (r5011);
    r4948 := (r4950 & r4952 & r4954 & r4956 & r4958 & r4960 & r4962 & r4964 & r4966 & r4968 & r4970 & r4972 & r4974 & r4976 & r4978 & r4980 & r4982 & r4984 & r4986 & r4988 & r4990 & r4992 & r4994 & r4996 & r4998 & r5000 & r5002 & r5004 & r5006 & r5008 & r5010 & r5012);
    return r4948;
  end rewire_MetaprogrammingRWw06ca6351_4947;
  function rewire_MetaprogrammingRWwd5a79147_4878 return std_logic_vector
  is
    variable r4943 : std_logic_vector(0 to 0) := (others => '0');
    variable r4942 : std_logic_vector(0 to 0) := (others => '0');
    variable r4941 : std_logic_vector(0 to 0) := (others => '0');
    variable r4940 : std_logic_vector(0 to 0) := (others => '0');
    variable r4939 : std_logic_vector(0 to 0) := (others => '0');
    variable r4938 : std_logic_vector(0 to 0) := (others => '0');
    variable r4937 : std_logic_vector(0 to 0) := (others => '0');
    variable r4936 : std_logic_vector(0 to 0) := (others => '0');
    variable r4935 : std_logic_vector(0 to 0) := (others => '0');
    variable r4934 : std_logic_vector(0 to 0) := (others => '0');
    variable r4933 : std_logic_vector(0 to 0) := (others => '0');
    variable r4932 : std_logic_vector(0 to 0) := (others => '0');
    variable r4931 : std_logic_vector(0 to 0) := (others => '0');
    variable r4930 : std_logic_vector(0 to 0) := (others => '0');
    variable r4929 : std_logic_vector(0 to 0) := (others => '0');
    variable r4928 : std_logic_vector(0 to 0) := (others => '0');
    variable r4927 : std_logic_vector(0 to 0) := (others => '0');
    variable r4926 : std_logic_vector(0 to 0) := (others => '0');
    variable r4925 : std_logic_vector(0 to 0) := (others => '0');
    variable r4924 : std_logic_vector(0 to 0) := (others => '0');
    variable r4923 : std_logic_vector(0 to 0) := (others => '0');
    variable r4922 : std_logic_vector(0 to 0) := (others => '0');
    variable r4921 : std_logic_vector(0 to 0) := (others => '0');
    variable r4920 : std_logic_vector(0 to 0) := (others => '0');
    variable r4919 : std_logic_vector(0 to 0) := (others => '0');
    variable r4918 : std_logic_vector(0 to 0) := (others => '0');
    variable r4917 : std_logic_vector(0 to 0) := (others => '0');
    variable r4916 : std_logic_vector(0 to 0) := (others => '0');
    variable r4915 : std_logic_vector(0 to 0) := (others => '0');
    variable r4914 : std_logic_vector(0 to 0) := (others => '0');
    variable r4913 : std_logic_vector(0 to 0) := (others => '0');
    variable r4912 : std_logic_vector(0 to 0) := (others => '0');
    variable r4911 : std_logic_vector(0 to 0) := (others => '0');
    variable r4910 : std_logic_vector(0 to 0) := (others => '0');
    variable r4909 : std_logic_vector(0 to 0) := (others => '0');
    variable r4908 : std_logic_vector(0 to 0) := (others => '0');
    variable r4907 : std_logic_vector(0 to 0) := (others => '0');
    variable r4906 : std_logic_vector(0 to 0) := (others => '0');
    variable r4905 : std_logic_vector(0 to 0) := (others => '0');
    variable r4904 : std_logic_vector(0 to 0) := (others => '0');
    variable r4903 : std_logic_vector(0 to 0) := (others => '0');
    variable r4902 : std_logic_vector(0 to 0) := (others => '0');
    variable r4901 : std_logic_vector(0 to 0) := (others => '0');
    variable r4900 : std_logic_vector(0 to 0) := (others => '0');
    variable r4899 : std_logic_vector(0 to 0) := (others => '0');
    variable r4898 : std_logic_vector(0 to 0) := (others => '0');
    variable r4897 : std_logic_vector(0 to 0) := (others => '0');
    variable r4896 : std_logic_vector(0 to 0) := (others => '0');
    variable r4895 : std_logic_vector(0 to 0) := (others => '0');
    variable r4894 : std_logic_vector(0 to 0) := (others => '0');
    variable r4893 : std_logic_vector(0 to 0) := (others => '0');
    variable r4892 : std_logic_vector(0 to 0) := (others => '0');
    variable r4891 : std_logic_vector(0 to 0) := (others => '0');
    variable r4890 : std_logic_vector(0 to 0) := (others => '0');
    variable r4889 : std_logic_vector(0 to 0) := (others => '0');
    variable r4888 : std_logic_vector(0 to 0) := (others => '0');
    variable r4887 : std_logic_vector(0 to 0) := (others => '0');
    variable r4886 : std_logic_vector(0 to 0) := (others => '0');
    variable r4885 : std_logic_vector(0 to 0) := (others => '0');
    variable r4884 : std_logic_vector(0 to 0) := (others => '0');
    variable r4883 : std_logic_vector(0 to 0) := (others => '0');
    variable r4882 : std_logic_vector(0 to 0) := (others => '0');
    variable r4881 : std_logic_vector(0 to 0) := (others => '0');
    variable r4880 : std_logic_vector(0 to 0) := (others => '0');
    variable r4879 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r4880 := "1";
    null;
    r4881 := (r4880);
    r4882 := "1";
    null;
    r4883 := (r4882);
    r4884 := "0";
    null;
    r4885 := (r4884);
    r4886 := "1";
    null;
    r4887 := (r4886);
    r4888 := "0";
    null;
    r4889 := (r4888);
    r4890 := "1";
    null;
    r4891 := (r4890);
    r4892 := "0";
    null;
    r4893 := (r4892);
    r4894 := "1";
    null;
    r4895 := (r4894);
    r4896 := "1";
    null;
    r4897 := (r4896);
    r4898 := "0";
    null;
    r4899 := (r4898);
    r4900 := "1";
    null;
    r4901 := (r4900);
    r4902 := "0";
    null;
    r4903 := (r4902);
    r4904 := "0";
    null;
    r4905 := (r4904);
    r4906 := "1";
    null;
    r4907 := (r4906);
    r4908 := "1";
    null;
    r4909 := (r4908);
    r4910 := "1";
    null;
    r4911 := (r4910);
    r4912 := "1";
    null;
    r4913 := (r4912);
    r4914 := "0";
    null;
    r4915 := (r4914);
    r4916 := "0";
    null;
    r4917 := (r4916);
    r4918 := "1";
    null;
    r4919 := (r4918);
    r4920 := "0";
    null;
    r4921 := (r4920);
    r4922 := "0";
    null;
    r4923 := (r4922);
    r4924 := "0";
    null;
    r4925 := (r4924);
    r4926 := "1";
    null;
    r4927 := (r4926);
    r4928 := "0";
    null;
    r4929 := (r4928);
    r4930 := "1";
    null;
    r4931 := (r4930);
    r4932 := "0";
    null;
    r4933 := (r4932);
    r4934 := "0";
    null;
    r4935 := (r4934);
    r4936 := "0";
    null;
    r4937 := (r4936);
    r4938 := "1";
    null;
    r4939 := (r4938);
    r4940 := "1";
    null;
    r4941 := (r4940);
    r4942 := "1";
    null;
    r4943 := (r4942);
    r4879 := (r4881 & r4883 & r4885 & r4887 & r4889 & r4891 & r4893 & r4895 & r4897 & r4899 & r4901 & r4903 & r4905 & r4907 & r4909 & r4911 & r4913 & r4915 & r4917 & r4919 & r4921 & r4923 & r4925 & r4927 & r4929 & r4931 & r4933 & r4935 & r4937 & r4939 & r4941 & r4943);
    return r4879;
  end rewire_MetaprogrammingRWwd5a79147_4878;
  function rewire_MetaprogrammingRWwc6e00bf3_4809 return std_logic_vector
  is
    variable r4874 : std_logic_vector(0 to 0) := (others => '0');
    variable r4873 : std_logic_vector(0 to 0) := (others => '0');
    variable r4872 : std_logic_vector(0 to 0) := (others => '0');
    variable r4871 : std_logic_vector(0 to 0) := (others => '0');
    variable r4870 : std_logic_vector(0 to 0) := (others => '0');
    variable r4869 : std_logic_vector(0 to 0) := (others => '0');
    variable r4868 : std_logic_vector(0 to 0) := (others => '0');
    variable r4867 : std_logic_vector(0 to 0) := (others => '0');
    variable r4866 : std_logic_vector(0 to 0) := (others => '0');
    variable r4865 : std_logic_vector(0 to 0) := (others => '0');
    variable r4864 : std_logic_vector(0 to 0) := (others => '0');
    variable r4863 : std_logic_vector(0 to 0) := (others => '0');
    variable r4862 : std_logic_vector(0 to 0) := (others => '0');
    variable r4861 : std_logic_vector(0 to 0) := (others => '0');
    variable r4860 : std_logic_vector(0 to 0) := (others => '0');
    variable r4859 : std_logic_vector(0 to 0) := (others => '0');
    variable r4858 : std_logic_vector(0 to 0) := (others => '0');
    variable r4857 : std_logic_vector(0 to 0) := (others => '0');
    variable r4856 : std_logic_vector(0 to 0) := (others => '0');
    variable r4855 : std_logic_vector(0 to 0) := (others => '0');
    variable r4854 : std_logic_vector(0 to 0) := (others => '0');
    variable r4853 : std_logic_vector(0 to 0) := (others => '0');
    variable r4852 : std_logic_vector(0 to 0) := (others => '0');
    variable r4851 : std_logic_vector(0 to 0) := (others => '0');
    variable r4850 : std_logic_vector(0 to 0) := (others => '0');
    variable r4849 : std_logic_vector(0 to 0) := (others => '0');
    variable r4848 : std_logic_vector(0 to 0) := (others => '0');
    variable r4847 : std_logic_vector(0 to 0) := (others => '0');
    variable r4846 : std_logic_vector(0 to 0) := (others => '0');
    variable r4845 : std_logic_vector(0 to 0) := (others => '0');
    variable r4844 : std_logic_vector(0 to 0) := (others => '0');
    variable r4843 : std_logic_vector(0 to 0) := (others => '0');
    variable r4842 : std_logic_vector(0 to 0) := (others => '0');
    variable r4841 : std_logic_vector(0 to 0) := (others => '0');
    variable r4840 : std_logic_vector(0 to 0) := (others => '0');
    variable r4839 : std_logic_vector(0 to 0) := (others => '0');
    variable r4838 : std_logic_vector(0 to 0) := (others => '0');
    variable r4837 : std_logic_vector(0 to 0) := (others => '0');
    variable r4836 : std_logic_vector(0 to 0) := (others => '0');
    variable r4835 : std_logic_vector(0 to 0) := (others => '0');
    variable r4834 : std_logic_vector(0 to 0) := (others => '0');
    variable r4833 : std_logic_vector(0 to 0) := (others => '0');
    variable r4832 : std_logic_vector(0 to 0) := (others => '0');
    variable r4831 : std_logic_vector(0 to 0) := (others => '0');
    variable r4830 : std_logic_vector(0 to 0) := (others => '0');
    variable r4829 : std_logic_vector(0 to 0) := (others => '0');
    variable r4828 : std_logic_vector(0 to 0) := (others => '0');
    variable r4827 : std_logic_vector(0 to 0) := (others => '0');
    variable r4826 : std_logic_vector(0 to 0) := (others => '0');
    variable r4825 : std_logic_vector(0 to 0) := (others => '0');
    variable r4824 : std_logic_vector(0 to 0) := (others => '0');
    variable r4823 : std_logic_vector(0 to 0) := (others => '0');
    variable r4822 : std_logic_vector(0 to 0) := (others => '0');
    variable r4821 : std_logic_vector(0 to 0) := (others => '0');
    variable r4820 : std_logic_vector(0 to 0) := (others => '0');
    variable r4819 : std_logic_vector(0 to 0) := (others => '0');
    variable r4818 : std_logic_vector(0 to 0) := (others => '0');
    variable r4817 : std_logic_vector(0 to 0) := (others => '0');
    variable r4816 : std_logic_vector(0 to 0) := (others => '0');
    variable r4815 : std_logic_vector(0 to 0) := (others => '0');
    variable r4814 : std_logic_vector(0 to 0) := (others => '0');
    variable r4813 : std_logic_vector(0 to 0) := (others => '0');
    variable r4812 : std_logic_vector(0 to 0) := (others => '0');
    variable r4811 : std_logic_vector(0 to 0) := (others => '0');
    variable r4810 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r4811 := "1";
    null;
    r4812 := (r4811);
    r4813 := "1";
    null;
    r4814 := (r4813);
    r4815 := "0";
    null;
    r4816 := (r4815);
    r4817 := "0";
    null;
    r4818 := (r4817);
    r4819 := "0";
    null;
    r4820 := (r4819);
    r4821 := "1";
    null;
    r4822 := (r4821);
    r4823 := "1";
    null;
    r4824 := (r4823);
    r4825 := "0";
    null;
    r4826 := (r4825);
    r4827 := "1";
    null;
    r4828 := (r4827);
    r4829 := "1";
    null;
    r4830 := (r4829);
    r4831 := "1";
    null;
    r4832 := (r4831);
    r4833 := "0";
    null;
    r4834 := (r4833);
    r4835 := "0";
    null;
    r4836 := (r4835);
    r4837 := "0";
    null;
    r4838 := (r4837);
    r4839 := "0";
    null;
    r4840 := (r4839);
    r4841 := "0";
    null;
    r4842 := (r4841);
    r4843 := "0";
    null;
    r4844 := (r4843);
    r4845 := "0";
    null;
    r4846 := (r4845);
    r4847 := "0";
    null;
    r4848 := (r4847);
    r4849 := "0";
    null;
    r4850 := (r4849);
    r4851 := "1";
    null;
    r4852 := (r4851);
    r4853 := "0";
    null;
    r4854 := (r4853);
    r4855 := "1";
    null;
    r4856 := (r4855);
    r4857 := "1";
    null;
    r4858 := (r4857);
    r4859 := "1";
    null;
    r4860 := (r4859);
    r4861 := "1";
    null;
    r4862 := (r4861);
    r4863 := "1";
    null;
    r4864 := (r4863);
    r4865 := "1";
    null;
    r4866 := (r4865);
    r4867 := "0";
    null;
    r4868 := (r4867);
    r4869 := "0";
    null;
    r4870 := (r4869);
    r4871 := "1";
    null;
    r4872 := (r4871);
    r4873 := "1";
    null;
    r4874 := (r4873);
    r4810 := (r4812 & r4814 & r4816 & r4818 & r4820 & r4822 & r4824 & r4826 & r4828 & r4830 & r4832 & r4834 & r4836 & r4838 & r4840 & r4842 & r4844 & r4846 & r4848 & r4850 & r4852 & r4854 & r4856 & r4858 & r4860 & r4862 & r4864 & r4866 & r4868 & r4870 & r4872 & r4874);
    return r4810;
  end rewire_MetaprogrammingRWwc6e00bf3_4809;
  function rewire_MetaprogrammingRWwbf597fc7_4740 return std_logic_vector
  is
    variable r4805 : std_logic_vector(0 to 0) := (others => '0');
    variable r4804 : std_logic_vector(0 to 0) := (others => '0');
    variable r4803 : std_logic_vector(0 to 0) := (others => '0');
    variable r4802 : std_logic_vector(0 to 0) := (others => '0');
    variable r4801 : std_logic_vector(0 to 0) := (others => '0');
    variable r4800 : std_logic_vector(0 to 0) := (others => '0');
    variable r4799 : std_logic_vector(0 to 0) := (others => '0');
    variable r4798 : std_logic_vector(0 to 0) := (others => '0');
    variable r4797 : std_logic_vector(0 to 0) := (others => '0');
    variable r4796 : std_logic_vector(0 to 0) := (others => '0');
    variable r4795 : std_logic_vector(0 to 0) := (others => '0');
    variable r4794 : std_logic_vector(0 to 0) := (others => '0');
    variable r4793 : std_logic_vector(0 to 0) := (others => '0');
    variable r4792 : std_logic_vector(0 to 0) := (others => '0');
    variable r4791 : std_logic_vector(0 to 0) := (others => '0');
    variable r4790 : std_logic_vector(0 to 0) := (others => '0');
    variable r4789 : std_logic_vector(0 to 0) := (others => '0');
    variable r4788 : std_logic_vector(0 to 0) := (others => '0');
    variable r4787 : std_logic_vector(0 to 0) := (others => '0');
    variable r4786 : std_logic_vector(0 to 0) := (others => '0');
    variable r4785 : std_logic_vector(0 to 0) := (others => '0');
    variable r4784 : std_logic_vector(0 to 0) := (others => '0');
    variable r4783 : std_logic_vector(0 to 0) := (others => '0');
    variable r4782 : std_logic_vector(0 to 0) := (others => '0');
    variable r4781 : std_logic_vector(0 to 0) := (others => '0');
    variable r4780 : std_logic_vector(0 to 0) := (others => '0');
    variable r4779 : std_logic_vector(0 to 0) := (others => '0');
    variable r4778 : std_logic_vector(0 to 0) := (others => '0');
    variable r4777 : std_logic_vector(0 to 0) := (others => '0');
    variable r4776 : std_logic_vector(0 to 0) := (others => '0');
    variable r4775 : std_logic_vector(0 to 0) := (others => '0');
    variable r4774 : std_logic_vector(0 to 0) := (others => '0');
    variable r4773 : std_logic_vector(0 to 0) := (others => '0');
    variable r4772 : std_logic_vector(0 to 0) := (others => '0');
    variable r4771 : std_logic_vector(0 to 0) := (others => '0');
    variable r4770 : std_logic_vector(0 to 0) := (others => '0');
    variable r4769 : std_logic_vector(0 to 0) := (others => '0');
    variable r4768 : std_logic_vector(0 to 0) := (others => '0');
    variable r4767 : std_logic_vector(0 to 0) := (others => '0');
    variable r4766 : std_logic_vector(0 to 0) := (others => '0');
    variable r4765 : std_logic_vector(0 to 0) := (others => '0');
    variable r4764 : std_logic_vector(0 to 0) := (others => '0');
    variable r4763 : std_logic_vector(0 to 0) := (others => '0');
    variable r4762 : std_logic_vector(0 to 0) := (others => '0');
    variable r4761 : std_logic_vector(0 to 0) := (others => '0');
    variable r4760 : std_logic_vector(0 to 0) := (others => '0');
    variable r4759 : std_logic_vector(0 to 0) := (others => '0');
    variable r4758 : std_logic_vector(0 to 0) := (others => '0');
    variable r4757 : std_logic_vector(0 to 0) := (others => '0');
    variable r4756 : std_logic_vector(0 to 0) := (others => '0');
    variable r4755 : std_logic_vector(0 to 0) := (others => '0');
    variable r4754 : std_logic_vector(0 to 0) := (others => '0');
    variable r4753 : std_logic_vector(0 to 0) := (others => '0');
    variable r4752 : std_logic_vector(0 to 0) := (others => '0');
    variable r4751 : std_logic_vector(0 to 0) := (others => '0');
    variable r4750 : std_logic_vector(0 to 0) := (others => '0');
    variable r4749 : std_logic_vector(0 to 0) := (others => '0');
    variable r4748 : std_logic_vector(0 to 0) := (others => '0');
    variable r4747 : std_logic_vector(0 to 0) := (others => '0');
    variable r4746 : std_logic_vector(0 to 0) := (others => '0');
    variable r4745 : std_logic_vector(0 to 0) := (others => '0');
    variable r4744 : std_logic_vector(0 to 0) := (others => '0');
    variable r4743 : std_logic_vector(0 to 0) := (others => '0');
    variable r4742 : std_logic_vector(0 to 0) := (others => '0');
    variable r4741 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r4742 := "1";
    null;
    r4743 := (r4742);
    r4744 := "0";
    null;
    r4745 := (r4744);
    r4746 := "1";
    null;
    r4747 := (r4746);
    r4748 := "1";
    null;
    r4749 := (r4748);
    r4750 := "1";
    null;
    r4751 := (r4750);
    r4752 := "1";
    null;
    r4753 := (r4752);
    r4754 := "1";
    null;
    r4755 := (r4754);
    r4756 := "1";
    null;
    r4757 := (r4756);
    r4758 := "0";
    null;
    r4759 := (r4758);
    r4760 := "1";
    null;
    r4761 := (r4760);
    r4762 := "0";
    null;
    r4763 := (r4762);
    r4764 := "1";
    null;
    r4765 := (r4764);
    r4766 := "1";
    null;
    r4767 := (r4766);
    r4768 := "0";
    null;
    r4769 := (r4768);
    r4770 := "0";
    null;
    r4771 := (r4770);
    r4772 := "1";
    null;
    r4773 := (r4772);
    r4774 := "0";
    null;
    r4775 := (r4774);
    r4776 := "1";
    null;
    r4777 := (r4776);
    r4778 := "1";
    null;
    r4779 := (r4778);
    r4780 := "1";
    null;
    r4781 := (r4780);
    r4782 := "1";
    null;
    r4783 := (r4782);
    r4784 := "1";
    null;
    r4785 := (r4784);
    r4786 := "1";
    null;
    r4787 := (r4786);
    r4788 := "1";
    null;
    r4789 := (r4788);
    r4790 := "1";
    null;
    r4791 := (r4790);
    r4792 := "1";
    null;
    r4793 := (r4792);
    r4794 := "0";
    null;
    r4795 := (r4794);
    r4796 := "0";
    null;
    r4797 := (r4796);
    r4798 := "0";
    null;
    r4799 := (r4798);
    r4800 := "1";
    null;
    r4801 := (r4800);
    r4802 := "1";
    null;
    r4803 := (r4802);
    r4804 := "1";
    null;
    r4805 := (r4804);
    r4741 := (r4743 & r4745 & r4747 & r4749 & r4751 & r4753 & r4755 & r4757 & r4759 & r4761 & r4763 & r4765 & r4767 & r4769 & r4771 & r4773 & r4775 & r4777 & r4779 & r4781 & r4783 & r4785 & r4787 & r4789 & r4791 & r4793 & r4795 & r4797 & r4799 & r4801 & r4803 & r4805);
    return r4741;
  end rewire_MetaprogrammingRWwbf597fc7_4740;
  function rewire_MetaprogrammingRWwb00327c8_4671 return std_logic_vector
  is
    variable r4736 : std_logic_vector(0 to 0) := (others => '0');
    variable r4735 : std_logic_vector(0 to 0) := (others => '0');
    variable r4734 : std_logic_vector(0 to 0) := (others => '0');
    variable r4733 : std_logic_vector(0 to 0) := (others => '0');
    variable r4732 : std_logic_vector(0 to 0) := (others => '0');
    variable r4731 : std_logic_vector(0 to 0) := (others => '0');
    variable r4730 : std_logic_vector(0 to 0) := (others => '0');
    variable r4729 : std_logic_vector(0 to 0) := (others => '0');
    variable r4728 : std_logic_vector(0 to 0) := (others => '0');
    variable r4727 : std_logic_vector(0 to 0) := (others => '0');
    variable r4726 : std_logic_vector(0 to 0) := (others => '0');
    variable r4725 : std_logic_vector(0 to 0) := (others => '0');
    variable r4724 : std_logic_vector(0 to 0) := (others => '0');
    variable r4723 : std_logic_vector(0 to 0) := (others => '0');
    variable r4722 : std_logic_vector(0 to 0) := (others => '0');
    variable r4721 : std_logic_vector(0 to 0) := (others => '0');
    variable r4720 : std_logic_vector(0 to 0) := (others => '0');
    variable r4719 : std_logic_vector(0 to 0) := (others => '0');
    variable r4718 : std_logic_vector(0 to 0) := (others => '0');
    variable r4717 : std_logic_vector(0 to 0) := (others => '0');
    variable r4716 : std_logic_vector(0 to 0) := (others => '0');
    variable r4715 : std_logic_vector(0 to 0) := (others => '0');
    variable r4714 : std_logic_vector(0 to 0) := (others => '0');
    variable r4713 : std_logic_vector(0 to 0) := (others => '0');
    variable r4712 : std_logic_vector(0 to 0) := (others => '0');
    variable r4711 : std_logic_vector(0 to 0) := (others => '0');
    variable r4710 : std_logic_vector(0 to 0) := (others => '0');
    variable r4709 : std_logic_vector(0 to 0) := (others => '0');
    variable r4708 : std_logic_vector(0 to 0) := (others => '0');
    variable r4707 : std_logic_vector(0 to 0) := (others => '0');
    variable r4706 : std_logic_vector(0 to 0) := (others => '0');
    variable r4705 : std_logic_vector(0 to 0) := (others => '0');
    variable r4704 : std_logic_vector(0 to 0) := (others => '0');
    variable r4703 : std_logic_vector(0 to 0) := (others => '0');
    variable r4702 : std_logic_vector(0 to 0) := (others => '0');
    variable r4701 : std_logic_vector(0 to 0) := (others => '0');
    variable r4700 : std_logic_vector(0 to 0) := (others => '0');
    variable r4699 : std_logic_vector(0 to 0) := (others => '0');
    variable r4698 : std_logic_vector(0 to 0) := (others => '0');
    variable r4697 : std_logic_vector(0 to 0) := (others => '0');
    variable r4696 : std_logic_vector(0 to 0) := (others => '0');
    variable r4695 : std_logic_vector(0 to 0) := (others => '0');
    variable r4694 : std_logic_vector(0 to 0) := (others => '0');
    variable r4693 : std_logic_vector(0 to 0) := (others => '0');
    variable r4692 : std_logic_vector(0 to 0) := (others => '0');
    variable r4691 : std_logic_vector(0 to 0) := (others => '0');
    variable r4690 : std_logic_vector(0 to 0) := (others => '0');
    variable r4689 : std_logic_vector(0 to 0) := (others => '0');
    variable r4688 : std_logic_vector(0 to 0) := (others => '0');
    variable r4687 : std_logic_vector(0 to 0) := (others => '0');
    variable r4686 : std_logic_vector(0 to 0) := (others => '0');
    variable r4685 : std_logic_vector(0 to 0) := (others => '0');
    variable r4684 : std_logic_vector(0 to 0) := (others => '0');
    variable r4683 : std_logic_vector(0 to 0) := (others => '0');
    variable r4682 : std_logic_vector(0 to 0) := (others => '0');
    variable r4681 : std_logic_vector(0 to 0) := (others => '0');
    variable r4680 : std_logic_vector(0 to 0) := (others => '0');
    variable r4679 : std_logic_vector(0 to 0) := (others => '0');
    variable r4678 : std_logic_vector(0 to 0) := (others => '0');
    variable r4677 : std_logic_vector(0 to 0) := (others => '0');
    variable r4676 : std_logic_vector(0 to 0) := (others => '0');
    variable r4675 : std_logic_vector(0 to 0) := (others => '0');
    variable r4674 : std_logic_vector(0 to 0) := (others => '0');
    variable r4673 : std_logic_vector(0 to 0) := (others => '0');
    variable r4672 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r4673 := "1";
    null;
    r4674 := (r4673);
    r4675 := "0";
    null;
    r4676 := (r4675);
    r4677 := "1";
    null;
    r4678 := (r4677);
    r4679 := "1";
    null;
    r4680 := (r4679);
    r4681 := "0";
    null;
    r4682 := (r4681);
    r4683 := "0";
    null;
    r4684 := (r4683);
    r4685 := "0";
    null;
    r4686 := (r4685);
    r4687 := "0";
    null;
    r4688 := (r4687);
    r4689 := "0";
    null;
    r4690 := (r4689);
    r4691 := "0";
    null;
    r4692 := (r4691);
    r4693 := "0";
    null;
    r4694 := (r4693);
    r4695 := "0";
    null;
    r4696 := (r4695);
    r4697 := "0";
    null;
    r4698 := (r4697);
    r4699 := "0";
    null;
    r4700 := (r4699);
    r4701 := "1";
    null;
    r4702 := (r4701);
    r4703 := "1";
    null;
    r4704 := (r4703);
    r4705 := "0";
    null;
    r4706 := (r4705);
    r4707 := "0";
    null;
    r4708 := (r4707);
    r4709 := "1";
    null;
    r4710 := (r4709);
    r4711 := "0";
    null;
    r4712 := (r4711);
    r4713 := "0";
    null;
    r4714 := (r4713);
    r4715 := "1";
    null;
    r4716 := (r4715);
    r4717 := "1";
    null;
    r4718 := (r4717);
    r4719 := "1";
    null;
    r4720 := (r4719);
    r4721 := "1";
    null;
    r4722 := (r4721);
    r4723 := "1";
    null;
    r4724 := (r4723);
    r4725 := "0";
    null;
    r4726 := (r4725);
    r4727 := "0";
    null;
    r4728 := (r4727);
    r4729 := "1";
    null;
    r4730 := (r4729);
    r4731 := "0";
    null;
    r4732 := (r4731);
    r4733 := "0";
    null;
    r4734 := (r4733);
    r4735 := "0";
    null;
    r4736 := (r4735);
    r4672 := (r4674 & r4676 & r4678 & r4680 & r4682 & r4684 & r4686 & r4688 & r4690 & r4692 & r4694 & r4696 & r4698 & r4700 & r4702 & r4704 & r4706 & r4708 & r4710 & r4712 & r4714 & r4716 & r4718 & r4720 & r4722 & r4724 & r4726 & r4728 & r4730 & r4732 & r4734 & r4736);
    return r4672;
  end rewire_MetaprogrammingRWwb00327c8_4671;
  function rewire_MetaprogrammingRWwa831c66d_4602 return std_logic_vector
  is
    variable r4667 : std_logic_vector(0 to 0) := (others => '0');
    variable r4666 : std_logic_vector(0 to 0) := (others => '0');
    variable r4665 : std_logic_vector(0 to 0) := (others => '0');
    variable r4664 : std_logic_vector(0 to 0) := (others => '0');
    variable r4663 : std_logic_vector(0 to 0) := (others => '0');
    variable r4662 : std_logic_vector(0 to 0) := (others => '0');
    variable r4661 : std_logic_vector(0 to 0) := (others => '0');
    variable r4660 : std_logic_vector(0 to 0) := (others => '0');
    variable r4659 : std_logic_vector(0 to 0) := (others => '0');
    variable r4658 : std_logic_vector(0 to 0) := (others => '0');
    variable r4657 : std_logic_vector(0 to 0) := (others => '0');
    variable r4656 : std_logic_vector(0 to 0) := (others => '0');
    variable r4655 : std_logic_vector(0 to 0) := (others => '0');
    variable r4654 : std_logic_vector(0 to 0) := (others => '0');
    variable r4653 : std_logic_vector(0 to 0) := (others => '0');
    variable r4652 : std_logic_vector(0 to 0) := (others => '0');
    variable r4651 : std_logic_vector(0 to 0) := (others => '0');
    variable r4650 : std_logic_vector(0 to 0) := (others => '0');
    variable r4649 : std_logic_vector(0 to 0) := (others => '0');
    variable r4648 : std_logic_vector(0 to 0) := (others => '0');
    variable r4647 : std_logic_vector(0 to 0) := (others => '0');
    variable r4646 : std_logic_vector(0 to 0) := (others => '0');
    variable r4645 : std_logic_vector(0 to 0) := (others => '0');
    variable r4644 : std_logic_vector(0 to 0) := (others => '0');
    variable r4643 : std_logic_vector(0 to 0) := (others => '0');
    variable r4642 : std_logic_vector(0 to 0) := (others => '0');
    variable r4641 : std_logic_vector(0 to 0) := (others => '0');
    variable r4640 : std_logic_vector(0 to 0) := (others => '0');
    variable r4639 : std_logic_vector(0 to 0) := (others => '0');
    variable r4638 : std_logic_vector(0 to 0) := (others => '0');
    variable r4637 : std_logic_vector(0 to 0) := (others => '0');
    variable r4636 : std_logic_vector(0 to 0) := (others => '0');
    variable r4635 : std_logic_vector(0 to 0) := (others => '0');
    variable r4634 : std_logic_vector(0 to 0) := (others => '0');
    variable r4633 : std_logic_vector(0 to 0) := (others => '0');
    variable r4632 : std_logic_vector(0 to 0) := (others => '0');
    variable r4631 : std_logic_vector(0 to 0) := (others => '0');
    variable r4630 : std_logic_vector(0 to 0) := (others => '0');
    variable r4629 : std_logic_vector(0 to 0) := (others => '0');
    variable r4628 : std_logic_vector(0 to 0) := (others => '0');
    variable r4627 : std_logic_vector(0 to 0) := (others => '0');
    variable r4626 : std_logic_vector(0 to 0) := (others => '0');
    variable r4625 : std_logic_vector(0 to 0) := (others => '0');
    variable r4624 : std_logic_vector(0 to 0) := (others => '0');
    variable r4623 : std_logic_vector(0 to 0) := (others => '0');
    variable r4622 : std_logic_vector(0 to 0) := (others => '0');
    variable r4621 : std_logic_vector(0 to 0) := (others => '0');
    variable r4620 : std_logic_vector(0 to 0) := (others => '0');
    variable r4619 : std_logic_vector(0 to 0) := (others => '0');
    variable r4618 : std_logic_vector(0 to 0) := (others => '0');
    variable r4617 : std_logic_vector(0 to 0) := (others => '0');
    variable r4616 : std_logic_vector(0 to 0) := (others => '0');
    variable r4615 : std_logic_vector(0 to 0) := (others => '0');
    variable r4614 : std_logic_vector(0 to 0) := (others => '0');
    variable r4613 : std_logic_vector(0 to 0) := (others => '0');
    variable r4612 : std_logic_vector(0 to 0) := (others => '0');
    variable r4611 : std_logic_vector(0 to 0) := (others => '0');
    variable r4610 : std_logic_vector(0 to 0) := (others => '0');
    variable r4609 : std_logic_vector(0 to 0) := (others => '0');
    variable r4608 : std_logic_vector(0 to 0) := (others => '0');
    variable r4607 : std_logic_vector(0 to 0) := (others => '0');
    variable r4606 : std_logic_vector(0 to 0) := (others => '0');
    variable r4605 : std_logic_vector(0 to 0) := (others => '0');
    variable r4604 : std_logic_vector(0 to 0) := (others => '0');
    variable r4603 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r4604 := "1";
    null;
    r4605 := (r4604);
    r4606 := "0";
    null;
    r4607 := (r4606);
    r4608 := "1";
    null;
    r4609 := (r4608);
    r4610 := "0";
    null;
    r4611 := (r4610);
    r4612 := "1";
    null;
    r4613 := (r4612);
    r4614 := "0";
    null;
    r4615 := (r4614);
    r4616 := "0";
    null;
    r4617 := (r4616);
    r4618 := "0";
    null;
    r4619 := (r4618);
    r4620 := "0";
    null;
    r4621 := (r4620);
    r4622 := "0";
    null;
    r4623 := (r4622);
    r4624 := "1";
    null;
    r4625 := (r4624);
    r4626 := "1";
    null;
    r4627 := (r4626);
    r4628 := "0";
    null;
    r4629 := (r4628);
    r4630 := "0";
    null;
    r4631 := (r4630);
    r4632 := "0";
    null;
    r4633 := (r4632);
    r4634 := "1";
    null;
    r4635 := (r4634);
    r4636 := "1";
    null;
    r4637 := (r4636);
    r4638 := "1";
    null;
    r4639 := (r4638);
    r4640 := "0";
    null;
    r4641 := (r4640);
    r4642 := "0";
    null;
    r4643 := (r4642);
    r4644 := "0";
    null;
    r4645 := (r4644);
    r4646 := "1";
    null;
    r4647 := (r4646);
    r4648 := "1";
    null;
    r4649 := (r4648);
    r4650 := "0";
    null;
    r4651 := (r4650);
    r4652 := "0";
    null;
    r4653 := (r4652);
    r4654 := "1";
    null;
    r4655 := (r4654);
    r4656 := "1";
    null;
    r4657 := (r4656);
    r4658 := "0";
    null;
    r4659 := (r4658);
    r4660 := "1";
    null;
    r4661 := (r4660);
    r4662 := "1";
    null;
    r4663 := (r4662);
    r4664 := "0";
    null;
    r4665 := (r4664);
    r4666 := "1";
    null;
    r4667 := (r4666);
    r4603 := (r4605 & r4607 & r4609 & r4611 & r4613 & r4615 & r4617 & r4619 & r4621 & r4623 & r4625 & r4627 & r4629 & r4631 & r4633 & r4635 & r4637 & r4639 & r4641 & r4643 & r4645 & r4647 & r4649 & r4651 & r4653 & r4655 & r4657 & r4659 & r4661 & r4663 & r4665 & r4667);
    return r4603;
  end rewire_MetaprogrammingRWwa831c66d_4602;
  function rewire_MetaprogrammingRWw983e5152_4533 return std_logic_vector
  is
    variable r4598 : std_logic_vector(0 to 0) := (others => '0');
    variable r4597 : std_logic_vector(0 to 0) := (others => '0');
    variable r4596 : std_logic_vector(0 to 0) := (others => '0');
    variable r4595 : std_logic_vector(0 to 0) := (others => '0');
    variable r4594 : std_logic_vector(0 to 0) := (others => '0');
    variable r4593 : std_logic_vector(0 to 0) := (others => '0');
    variable r4592 : std_logic_vector(0 to 0) := (others => '0');
    variable r4591 : std_logic_vector(0 to 0) := (others => '0');
    variable r4590 : std_logic_vector(0 to 0) := (others => '0');
    variable r4589 : std_logic_vector(0 to 0) := (others => '0');
    variable r4588 : std_logic_vector(0 to 0) := (others => '0');
    variable r4587 : std_logic_vector(0 to 0) := (others => '0');
    variable r4586 : std_logic_vector(0 to 0) := (others => '0');
    variable r4585 : std_logic_vector(0 to 0) := (others => '0');
    variable r4584 : std_logic_vector(0 to 0) := (others => '0');
    variable r4583 : std_logic_vector(0 to 0) := (others => '0');
    variable r4582 : std_logic_vector(0 to 0) := (others => '0');
    variable r4581 : std_logic_vector(0 to 0) := (others => '0');
    variable r4580 : std_logic_vector(0 to 0) := (others => '0');
    variable r4579 : std_logic_vector(0 to 0) := (others => '0');
    variable r4578 : std_logic_vector(0 to 0) := (others => '0');
    variable r4577 : std_logic_vector(0 to 0) := (others => '0');
    variable r4576 : std_logic_vector(0 to 0) := (others => '0');
    variable r4575 : std_logic_vector(0 to 0) := (others => '0');
    variable r4574 : std_logic_vector(0 to 0) := (others => '0');
    variable r4573 : std_logic_vector(0 to 0) := (others => '0');
    variable r4572 : std_logic_vector(0 to 0) := (others => '0');
    variable r4571 : std_logic_vector(0 to 0) := (others => '0');
    variable r4570 : std_logic_vector(0 to 0) := (others => '0');
    variable r4569 : std_logic_vector(0 to 0) := (others => '0');
    variable r4568 : std_logic_vector(0 to 0) := (others => '0');
    variable r4567 : std_logic_vector(0 to 0) := (others => '0');
    variable r4566 : std_logic_vector(0 to 0) := (others => '0');
    variable r4565 : std_logic_vector(0 to 0) := (others => '0');
    variable r4564 : std_logic_vector(0 to 0) := (others => '0');
    variable r4563 : std_logic_vector(0 to 0) := (others => '0');
    variable r4562 : std_logic_vector(0 to 0) := (others => '0');
    variable r4561 : std_logic_vector(0 to 0) := (others => '0');
    variable r4560 : std_logic_vector(0 to 0) := (others => '0');
    variable r4559 : std_logic_vector(0 to 0) := (others => '0');
    variable r4558 : std_logic_vector(0 to 0) := (others => '0');
    variable r4557 : std_logic_vector(0 to 0) := (others => '0');
    variable r4556 : std_logic_vector(0 to 0) := (others => '0');
    variable r4555 : std_logic_vector(0 to 0) := (others => '0');
    variable r4554 : std_logic_vector(0 to 0) := (others => '0');
    variable r4553 : std_logic_vector(0 to 0) := (others => '0');
    variable r4552 : std_logic_vector(0 to 0) := (others => '0');
    variable r4551 : std_logic_vector(0 to 0) := (others => '0');
    variable r4550 : std_logic_vector(0 to 0) := (others => '0');
    variable r4549 : std_logic_vector(0 to 0) := (others => '0');
    variable r4548 : std_logic_vector(0 to 0) := (others => '0');
    variable r4547 : std_logic_vector(0 to 0) := (others => '0');
    variable r4546 : std_logic_vector(0 to 0) := (others => '0');
    variable r4545 : std_logic_vector(0 to 0) := (others => '0');
    variable r4544 : std_logic_vector(0 to 0) := (others => '0');
    variable r4543 : std_logic_vector(0 to 0) := (others => '0');
    variable r4542 : std_logic_vector(0 to 0) := (others => '0');
    variable r4541 : std_logic_vector(0 to 0) := (others => '0');
    variable r4540 : std_logic_vector(0 to 0) := (others => '0');
    variable r4539 : std_logic_vector(0 to 0) := (others => '0');
    variable r4538 : std_logic_vector(0 to 0) := (others => '0');
    variable r4537 : std_logic_vector(0 to 0) := (others => '0');
    variable r4536 : std_logic_vector(0 to 0) := (others => '0');
    variable r4535 : std_logic_vector(0 to 0) := (others => '0');
    variable r4534 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r4535 := "1";
    null;
    r4536 := (r4535);
    r4537 := "0";
    null;
    r4538 := (r4537);
    r4539 := "0";
    null;
    r4540 := (r4539);
    r4541 := "1";
    null;
    r4542 := (r4541);
    r4543 := "1";
    null;
    r4544 := (r4543);
    r4545 := "0";
    null;
    r4546 := (r4545);
    r4547 := "0";
    null;
    r4548 := (r4547);
    r4549 := "0";
    null;
    r4550 := (r4549);
    r4551 := "0";
    null;
    r4552 := (r4551);
    r4553 := "0";
    null;
    r4554 := (r4553);
    r4555 := "1";
    null;
    r4556 := (r4555);
    r4557 := "1";
    null;
    r4558 := (r4557);
    r4559 := "1";
    null;
    r4560 := (r4559);
    r4561 := "1";
    null;
    r4562 := (r4561);
    r4563 := "1";
    null;
    r4564 := (r4563);
    r4565 := "0";
    null;
    r4566 := (r4565);
    r4567 := "0";
    null;
    r4568 := (r4567);
    r4569 := "1";
    null;
    r4570 := (r4569);
    r4571 := "0";
    null;
    r4572 := (r4571);
    r4573 := "1";
    null;
    r4574 := (r4573);
    r4575 := "0";
    null;
    r4576 := (r4575);
    r4577 := "0";
    null;
    r4578 := (r4577);
    r4579 := "0";
    null;
    r4580 := (r4579);
    r4581 := "1";
    null;
    r4582 := (r4581);
    r4583 := "0";
    null;
    r4584 := (r4583);
    r4585 := "1";
    null;
    r4586 := (r4585);
    r4587 := "0";
    null;
    r4588 := (r4587);
    r4589 := "1";
    null;
    r4590 := (r4589);
    r4591 := "0";
    null;
    r4592 := (r4591);
    r4593 := "0";
    null;
    r4594 := (r4593);
    r4595 := "1";
    null;
    r4596 := (r4595);
    r4597 := "0";
    null;
    r4598 := (r4597);
    r4534 := (r4536 & r4538 & r4540 & r4542 & r4544 & r4546 & r4548 & r4550 & r4552 & r4554 & r4556 & r4558 & r4560 & r4562 & r4564 & r4566 & r4568 & r4570 & r4572 & r4574 & r4576 & r4578 & r4580 & r4582 & r4584 & r4586 & r4588 & r4590 & r4592 & r4594 & r4596 & r4598);
    return r4534;
  end rewire_MetaprogrammingRWw983e5152_4533;
  function rewire_MetaprogrammingRWw76f988da_4464 return std_logic_vector
  is
    variable r4529 : std_logic_vector(0 to 0) := (others => '0');
    variable r4528 : std_logic_vector(0 to 0) := (others => '0');
    variable r4527 : std_logic_vector(0 to 0) := (others => '0');
    variable r4526 : std_logic_vector(0 to 0) := (others => '0');
    variable r4525 : std_logic_vector(0 to 0) := (others => '0');
    variable r4524 : std_logic_vector(0 to 0) := (others => '0');
    variable r4523 : std_logic_vector(0 to 0) := (others => '0');
    variable r4522 : std_logic_vector(0 to 0) := (others => '0');
    variable r4521 : std_logic_vector(0 to 0) := (others => '0');
    variable r4520 : std_logic_vector(0 to 0) := (others => '0');
    variable r4519 : std_logic_vector(0 to 0) := (others => '0');
    variable r4518 : std_logic_vector(0 to 0) := (others => '0');
    variable r4517 : std_logic_vector(0 to 0) := (others => '0');
    variable r4516 : std_logic_vector(0 to 0) := (others => '0');
    variable r4515 : std_logic_vector(0 to 0) := (others => '0');
    variable r4514 : std_logic_vector(0 to 0) := (others => '0');
    variable r4513 : std_logic_vector(0 to 0) := (others => '0');
    variable r4512 : std_logic_vector(0 to 0) := (others => '0');
    variable r4511 : std_logic_vector(0 to 0) := (others => '0');
    variable r4510 : std_logic_vector(0 to 0) := (others => '0');
    variable r4509 : std_logic_vector(0 to 0) := (others => '0');
    variable r4508 : std_logic_vector(0 to 0) := (others => '0');
    variable r4507 : std_logic_vector(0 to 0) := (others => '0');
    variable r4506 : std_logic_vector(0 to 0) := (others => '0');
    variable r4505 : std_logic_vector(0 to 0) := (others => '0');
    variable r4504 : std_logic_vector(0 to 0) := (others => '0');
    variable r4503 : std_logic_vector(0 to 0) := (others => '0');
    variable r4502 : std_logic_vector(0 to 0) := (others => '0');
    variable r4501 : std_logic_vector(0 to 0) := (others => '0');
    variable r4500 : std_logic_vector(0 to 0) := (others => '0');
    variable r4499 : std_logic_vector(0 to 0) := (others => '0');
    variable r4498 : std_logic_vector(0 to 0) := (others => '0');
    variable r4497 : std_logic_vector(0 to 0) := (others => '0');
    variable r4496 : std_logic_vector(0 to 0) := (others => '0');
    variable r4495 : std_logic_vector(0 to 0) := (others => '0');
    variable r4494 : std_logic_vector(0 to 0) := (others => '0');
    variable r4493 : std_logic_vector(0 to 0) := (others => '0');
    variable r4492 : std_logic_vector(0 to 0) := (others => '0');
    variable r4491 : std_logic_vector(0 to 0) := (others => '0');
    variable r4490 : std_logic_vector(0 to 0) := (others => '0');
    variable r4489 : std_logic_vector(0 to 0) := (others => '0');
    variable r4488 : std_logic_vector(0 to 0) := (others => '0');
    variable r4487 : std_logic_vector(0 to 0) := (others => '0');
    variable r4486 : std_logic_vector(0 to 0) := (others => '0');
    variable r4485 : std_logic_vector(0 to 0) := (others => '0');
    variable r4484 : std_logic_vector(0 to 0) := (others => '0');
    variable r4483 : std_logic_vector(0 to 0) := (others => '0');
    variable r4482 : std_logic_vector(0 to 0) := (others => '0');
    variable r4481 : std_logic_vector(0 to 0) := (others => '0');
    variable r4480 : std_logic_vector(0 to 0) := (others => '0');
    variable r4479 : std_logic_vector(0 to 0) := (others => '0');
    variable r4478 : std_logic_vector(0 to 0) := (others => '0');
    variable r4477 : std_logic_vector(0 to 0) := (others => '0');
    variable r4476 : std_logic_vector(0 to 0) := (others => '0');
    variable r4475 : std_logic_vector(0 to 0) := (others => '0');
    variable r4474 : std_logic_vector(0 to 0) := (others => '0');
    variable r4473 : std_logic_vector(0 to 0) := (others => '0');
    variable r4472 : std_logic_vector(0 to 0) := (others => '0');
    variable r4471 : std_logic_vector(0 to 0) := (others => '0');
    variable r4470 : std_logic_vector(0 to 0) := (others => '0');
    variable r4469 : std_logic_vector(0 to 0) := (others => '0');
    variable r4468 : std_logic_vector(0 to 0) := (others => '0');
    variable r4467 : std_logic_vector(0 to 0) := (others => '0');
    variable r4466 : std_logic_vector(0 to 0) := (others => '0');
    variable r4465 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r4466 := "0";
    null;
    r4467 := (r4466);
    r4468 := "1";
    null;
    r4469 := (r4468);
    r4470 := "1";
    null;
    r4471 := (r4470);
    r4472 := "1";
    null;
    r4473 := (r4472);
    r4474 := "0";
    null;
    r4475 := (r4474);
    r4476 := "1";
    null;
    r4477 := (r4476);
    r4478 := "1";
    null;
    r4479 := (r4478);
    r4480 := "0";
    null;
    r4481 := (r4480);
    r4482 := "1";
    null;
    r4483 := (r4482);
    r4484 := "1";
    null;
    r4485 := (r4484);
    r4486 := "1";
    null;
    r4487 := (r4486);
    r4488 := "1";
    null;
    r4489 := (r4488);
    r4490 := "1";
    null;
    r4491 := (r4490);
    r4492 := "0";
    null;
    r4493 := (r4492);
    r4494 := "0";
    null;
    r4495 := (r4494);
    r4496 := "1";
    null;
    r4497 := (r4496);
    r4498 := "1";
    null;
    r4499 := (r4498);
    r4500 := "0";
    null;
    r4501 := (r4500);
    r4502 := "0";
    null;
    r4503 := (r4502);
    r4504 := "0";
    null;
    r4505 := (r4504);
    r4506 := "1";
    null;
    r4507 := (r4506);
    r4508 := "0";
    null;
    r4509 := (r4508);
    r4510 := "0";
    null;
    r4511 := (r4510);
    r4512 := "0";
    null;
    r4513 := (r4512);
    r4514 := "1";
    null;
    r4515 := (r4514);
    r4516 := "1";
    null;
    r4517 := (r4516);
    r4518 := "0";
    null;
    r4519 := (r4518);
    r4520 := "1";
    null;
    r4521 := (r4520);
    r4522 := "1";
    null;
    r4523 := (r4522);
    r4524 := "0";
    null;
    r4525 := (r4524);
    r4526 := "1";
    null;
    r4527 := (r4526);
    r4528 := "0";
    null;
    r4529 := (r4528);
    r4465 := (r4467 & r4469 & r4471 & r4473 & r4475 & r4477 & r4479 & r4481 & r4483 & r4485 & r4487 & r4489 & r4491 & r4493 & r4495 & r4497 & r4499 & r4501 & r4503 & r4505 & r4507 & r4509 & r4511 & r4513 & r4515 & r4517 & r4519 & r4521 & r4523 & r4525 & r4527 & r4529);
    return r4465;
  end rewire_MetaprogrammingRWw76f988da_4464;
  function rewire_MetaprogrammingRWw5cb0a9dc_4395 return std_logic_vector
  is
    variable r4460 : std_logic_vector(0 to 0) := (others => '0');
    variable r4459 : std_logic_vector(0 to 0) := (others => '0');
    variable r4458 : std_logic_vector(0 to 0) := (others => '0');
    variable r4457 : std_logic_vector(0 to 0) := (others => '0');
    variable r4456 : std_logic_vector(0 to 0) := (others => '0');
    variable r4455 : std_logic_vector(0 to 0) := (others => '0');
    variable r4454 : std_logic_vector(0 to 0) := (others => '0');
    variable r4453 : std_logic_vector(0 to 0) := (others => '0');
    variable r4452 : std_logic_vector(0 to 0) := (others => '0');
    variable r4451 : std_logic_vector(0 to 0) := (others => '0');
    variable r4450 : std_logic_vector(0 to 0) := (others => '0');
    variable r4449 : std_logic_vector(0 to 0) := (others => '0');
    variable r4448 : std_logic_vector(0 to 0) := (others => '0');
    variable r4447 : std_logic_vector(0 to 0) := (others => '0');
    variable r4446 : std_logic_vector(0 to 0) := (others => '0');
    variable r4445 : std_logic_vector(0 to 0) := (others => '0');
    variable r4444 : std_logic_vector(0 to 0) := (others => '0');
    variable r4443 : std_logic_vector(0 to 0) := (others => '0');
    variable r4442 : std_logic_vector(0 to 0) := (others => '0');
    variable r4441 : std_logic_vector(0 to 0) := (others => '0');
    variable r4440 : std_logic_vector(0 to 0) := (others => '0');
    variable r4439 : std_logic_vector(0 to 0) := (others => '0');
    variable r4438 : std_logic_vector(0 to 0) := (others => '0');
    variable r4437 : std_logic_vector(0 to 0) := (others => '0');
    variable r4436 : std_logic_vector(0 to 0) := (others => '0');
    variable r4435 : std_logic_vector(0 to 0) := (others => '0');
    variable r4434 : std_logic_vector(0 to 0) := (others => '0');
    variable r4433 : std_logic_vector(0 to 0) := (others => '0');
    variable r4432 : std_logic_vector(0 to 0) := (others => '0');
    variable r4431 : std_logic_vector(0 to 0) := (others => '0');
    variable r4430 : std_logic_vector(0 to 0) := (others => '0');
    variable r4429 : std_logic_vector(0 to 0) := (others => '0');
    variable r4428 : std_logic_vector(0 to 0) := (others => '0');
    variable r4427 : std_logic_vector(0 to 0) := (others => '0');
    variable r4426 : std_logic_vector(0 to 0) := (others => '0');
    variable r4425 : std_logic_vector(0 to 0) := (others => '0');
    variable r4424 : std_logic_vector(0 to 0) := (others => '0');
    variable r4423 : std_logic_vector(0 to 0) := (others => '0');
    variable r4422 : std_logic_vector(0 to 0) := (others => '0');
    variable r4421 : std_logic_vector(0 to 0) := (others => '0');
    variable r4420 : std_logic_vector(0 to 0) := (others => '0');
    variable r4419 : std_logic_vector(0 to 0) := (others => '0');
    variable r4418 : std_logic_vector(0 to 0) := (others => '0');
    variable r4417 : std_logic_vector(0 to 0) := (others => '0');
    variable r4416 : std_logic_vector(0 to 0) := (others => '0');
    variable r4415 : std_logic_vector(0 to 0) := (others => '0');
    variable r4414 : std_logic_vector(0 to 0) := (others => '0');
    variable r4413 : std_logic_vector(0 to 0) := (others => '0');
    variable r4412 : std_logic_vector(0 to 0) := (others => '0');
    variable r4411 : std_logic_vector(0 to 0) := (others => '0');
    variable r4410 : std_logic_vector(0 to 0) := (others => '0');
    variable r4409 : std_logic_vector(0 to 0) := (others => '0');
    variable r4408 : std_logic_vector(0 to 0) := (others => '0');
    variable r4407 : std_logic_vector(0 to 0) := (others => '0');
    variable r4406 : std_logic_vector(0 to 0) := (others => '0');
    variable r4405 : std_logic_vector(0 to 0) := (others => '0');
    variable r4404 : std_logic_vector(0 to 0) := (others => '0');
    variable r4403 : std_logic_vector(0 to 0) := (others => '0');
    variable r4402 : std_logic_vector(0 to 0) := (others => '0');
    variable r4401 : std_logic_vector(0 to 0) := (others => '0');
    variable r4400 : std_logic_vector(0 to 0) := (others => '0');
    variable r4399 : std_logic_vector(0 to 0) := (others => '0');
    variable r4398 : std_logic_vector(0 to 0) := (others => '0');
    variable r4397 : std_logic_vector(0 to 0) := (others => '0');
    variable r4396 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r4397 := "0";
    null;
    r4398 := (r4397);
    r4399 := "1";
    null;
    r4400 := (r4399);
    r4401 := "0";
    null;
    r4402 := (r4401);
    r4403 := "1";
    null;
    r4404 := (r4403);
    r4405 := "1";
    null;
    r4406 := (r4405);
    r4407 := "1";
    null;
    r4408 := (r4407);
    r4409 := "0";
    null;
    r4410 := (r4409);
    r4411 := "0";
    null;
    r4412 := (r4411);
    r4413 := "1";
    null;
    r4414 := (r4413);
    r4415 := "0";
    null;
    r4416 := (r4415);
    r4417 := "1";
    null;
    r4418 := (r4417);
    r4419 := "1";
    null;
    r4420 := (r4419);
    r4421 := "0";
    null;
    r4422 := (r4421);
    r4423 := "0";
    null;
    r4424 := (r4423);
    r4425 := "0";
    null;
    r4426 := (r4425);
    r4427 := "0";
    null;
    r4428 := (r4427);
    r4429 := "1";
    null;
    r4430 := (r4429);
    r4431 := "0";
    null;
    r4432 := (r4431);
    r4433 := "1";
    null;
    r4434 := (r4433);
    r4435 := "0";
    null;
    r4436 := (r4435);
    r4437 := "1";
    null;
    r4438 := (r4437);
    r4439 := "0";
    null;
    r4440 := (r4439);
    r4441 := "0";
    null;
    r4442 := (r4441);
    r4443 := "1";
    null;
    r4444 := (r4443);
    r4445 := "1";
    null;
    r4446 := (r4445);
    r4447 := "1";
    null;
    r4448 := (r4447);
    r4449 := "0";
    null;
    r4450 := (r4449);
    r4451 := "1";
    null;
    r4452 := (r4451);
    r4453 := "1";
    null;
    r4454 := (r4453);
    r4455 := "1";
    null;
    r4456 := (r4455);
    r4457 := "0";
    null;
    r4458 := (r4457);
    r4459 := "0";
    null;
    r4460 := (r4459);
    r4396 := (r4398 & r4400 & r4402 & r4404 & r4406 & r4408 & r4410 & r4412 & r4414 & r4416 & r4418 & r4420 & r4422 & r4424 & r4426 & r4428 & r4430 & r4432 & r4434 & r4436 & r4438 & r4440 & r4442 & r4444 & r4446 & r4448 & r4450 & r4452 & r4454 & r4456 & r4458 & r4460);
    return r4396;
  end rewire_MetaprogrammingRWw5cb0a9dc_4395;
  function rewire_MetaprogrammingRWw4a7484aa_4326 return std_logic_vector
  is
    variable r4391 : std_logic_vector(0 to 0) := (others => '0');
    variable r4390 : std_logic_vector(0 to 0) := (others => '0');
    variable r4389 : std_logic_vector(0 to 0) := (others => '0');
    variable r4388 : std_logic_vector(0 to 0) := (others => '0');
    variable r4387 : std_logic_vector(0 to 0) := (others => '0');
    variable r4386 : std_logic_vector(0 to 0) := (others => '0');
    variable r4385 : std_logic_vector(0 to 0) := (others => '0');
    variable r4384 : std_logic_vector(0 to 0) := (others => '0');
    variable r4383 : std_logic_vector(0 to 0) := (others => '0');
    variable r4382 : std_logic_vector(0 to 0) := (others => '0');
    variable r4381 : std_logic_vector(0 to 0) := (others => '0');
    variable r4380 : std_logic_vector(0 to 0) := (others => '0');
    variable r4379 : std_logic_vector(0 to 0) := (others => '0');
    variable r4378 : std_logic_vector(0 to 0) := (others => '0');
    variable r4377 : std_logic_vector(0 to 0) := (others => '0');
    variable r4376 : std_logic_vector(0 to 0) := (others => '0');
    variable r4375 : std_logic_vector(0 to 0) := (others => '0');
    variable r4374 : std_logic_vector(0 to 0) := (others => '0');
    variable r4373 : std_logic_vector(0 to 0) := (others => '0');
    variable r4372 : std_logic_vector(0 to 0) := (others => '0');
    variable r4371 : std_logic_vector(0 to 0) := (others => '0');
    variable r4370 : std_logic_vector(0 to 0) := (others => '0');
    variable r4369 : std_logic_vector(0 to 0) := (others => '0');
    variable r4368 : std_logic_vector(0 to 0) := (others => '0');
    variable r4367 : std_logic_vector(0 to 0) := (others => '0');
    variable r4366 : std_logic_vector(0 to 0) := (others => '0');
    variable r4365 : std_logic_vector(0 to 0) := (others => '0');
    variable r4364 : std_logic_vector(0 to 0) := (others => '0');
    variable r4363 : std_logic_vector(0 to 0) := (others => '0');
    variable r4362 : std_logic_vector(0 to 0) := (others => '0');
    variable r4361 : std_logic_vector(0 to 0) := (others => '0');
    variable r4360 : std_logic_vector(0 to 0) := (others => '0');
    variable r4359 : std_logic_vector(0 to 0) := (others => '0');
    variable r4358 : std_logic_vector(0 to 0) := (others => '0');
    variable r4357 : std_logic_vector(0 to 0) := (others => '0');
    variable r4356 : std_logic_vector(0 to 0) := (others => '0');
    variable r4355 : std_logic_vector(0 to 0) := (others => '0');
    variable r4354 : std_logic_vector(0 to 0) := (others => '0');
    variable r4353 : std_logic_vector(0 to 0) := (others => '0');
    variable r4352 : std_logic_vector(0 to 0) := (others => '0');
    variable r4351 : std_logic_vector(0 to 0) := (others => '0');
    variable r4350 : std_logic_vector(0 to 0) := (others => '0');
    variable r4349 : std_logic_vector(0 to 0) := (others => '0');
    variable r4348 : std_logic_vector(0 to 0) := (others => '0');
    variable r4347 : std_logic_vector(0 to 0) := (others => '0');
    variable r4346 : std_logic_vector(0 to 0) := (others => '0');
    variable r4345 : std_logic_vector(0 to 0) := (others => '0');
    variable r4344 : std_logic_vector(0 to 0) := (others => '0');
    variable r4343 : std_logic_vector(0 to 0) := (others => '0');
    variable r4342 : std_logic_vector(0 to 0) := (others => '0');
    variable r4341 : std_logic_vector(0 to 0) := (others => '0');
    variable r4340 : std_logic_vector(0 to 0) := (others => '0');
    variable r4339 : std_logic_vector(0 to 0) := (others => '0');
    variable r4338 : std_logic_vector(0 to 0) := (others => '0');
    variable r4337 : std_logic_vector(0 to 0) := (others => '0');
    variable r4336 : std_logic_vector(0 to 0) := (others => '0');
    variable r4335 : std_logic_vector(0 to 0) := (others => '0');
    variable r4334 : std_logic_vector(0 to 0) := (others => '0');
    variable r4333 : std_logic_vector(0 to 0) := (others => '0');
    variable r4332 : std_logic_vector(0 to 0) := (others => '0');
    variable r4331 : std_logic_vector(0 to 0) := (others => '0');
    variable r4330 : std_logic_vector(0 to 0) := (others => '0');
    variable r4329 : std_logic_vector(0 to 0) := (others => '0');
    variable r4328 : std_logic_vector(0 to 0) := (others => '0');
    variable r4327 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r4328 := "0";
    null;
    r4329 := (r4328);
    r4330 := "1";
    null;
    r4331 := (r4330);
    r4332 := "0";
    null;
    r4333 := (r4332);
    r4334 := "0";
    null;
    r4335 := (r4334);
    r4336 := "1";
    null;
    r4337 := (r4336);
    r4338 := "0";
    null;
    r4339 := (r4338);
    r4340 := "1";
    null;
    r4341 := (r4340);
    r4342 := "0";
    null;
    r4343 := (r4342);
    r4344 := "0";
    null;
    r4345 := (r4344);
    r4346 := "1";
    null;
    r4347 := (r4346);
    r4348 := "1";
    null;
    r4349 := (r4348);
    r4350 := "1";
    null;
    r4351 := (r4350);
    r4352 := "0";
    null;
    r4353 := (r4352);
    r4354 := "1";
    null;
    r4355 := (r4354);
    r4356 := "0";
    null;
    r4357 := (r4356);
    r4358 := "0";
    null;
    r4359 := (r4358);
    r4360 := "1";
    null;
    r4361 := (r4360);
    r4362 := "0";
    null;
    r4363 := (r4362);
    r4364 := "0";
    null;
    r4365 := (r4364);
    r4366 := "0";
    null;
    r4367 := (r4366);
    r4368 := "0";
    null;
    r4369 := (r4368);
    r4370 := "1";
    null;
    r4371 := (r4370);
    r4372 := "0";
    null;
    r4373 := (r4372);
    r4374 := "0";
    null;
    r4375 := (r4374);
    r4376 := "1";
    null;
    r4377 := (r4376);
    r4378 := "0";
    null;
    r4379 := (r4378);
    r4380 := "1";
    null;
    r4381 := (r4380);
    r4382 := "0";
    null;
    r4383 := (r4382);
    r4384 := "1";
    null;
    r4385 := (r4384);
    r4386 := "0";
    null;
    r4387 := (r4386);
    r4388 := "1";
    null;
    r4389 := (r4388);
    r4390 := "0";
    null;
    r4391 := (r4390);
    r4327 := (r4329 & r4331 & r4333 & r4335 & r4337 & r4339 & r4341 & r4343 & r4345 & r4347 & r4349 & r4351 & r4353 & r4355 & r4357 & r4359 & r4361 & r4363 & r4365 & r4367 & r4369 & r4371 & r4373 & r4375 & r4377 & r4379 & r4381 & r4383 & r4385 & r4387 & r4389 & r4391);
    return r4327;
  end rewire_MetaprogrammingRWw4a7484aa_4326;
  function rewire_MetaprogrammingRWw2de92c6f_4257 return std_logic_vector
  is
    variable r4322 : std_logic_vector(0 to 0) := (others => '0');
    variable r4321 : std_logic_vector(0 to 0) := (others => '0');
    variable r4320 : std_logic_vector(0 to 0) := (others => '0');
    variable r4319 : std_logic_vector(0 to 0) := (others => '0');
    variable r4318 : std_logic_vector(0 to 0) := (others => '0');
    variable r4317 : std_logic_vector(0 to 0) := (others => '0');
    variable r4316 : std_logic_vector(0 to 0) := (others => '0');
    variable r4315 : std_logic_vector(0 to 0) := (others => '0');
    variable r4314 : std_logic_vector(0 to 0) := (others => '0');
    variable r4313 : std_logic_vector(0 to 0) := (others => '0');
    variable r4312 : std_logic_vector(0 to 0) := (others => '0');
    variable r4311 : std_logic_vector(0 to 0) := (others => '0');
    variable r4310 : std_logic_vector(0 to 0) := (others => '0');
    variable r4309 : std_logic_vector(0 to 0) := (others => '0');
    variable r4308 : std_logic_vector(0 to 0) := (others => '0');
    variable r4307 : std_logic_vector(0 to 0) := (others => '0');
    variable r4306 : std_logic_vector(0 to 0) := (others => '0');
    variable r4305 : std_logic_vector(0 to 0) := (others => '0');
    variable r4304 : std_logic_vector(0 to 0) := (others => '0');
    variable r4303 : std_logic_vector(0 to 0) := (others => '0');
    variable r4302 : std_logic_vector(0 to 0) := (others => '0');
    variable r4301 : std_logic_vector(0 to 0) := (others => '0');
    variable r4300 : std_logic_vector(0 to 0) := (others => '0');
    variable r4299 : std_logic_vector(0 to 0) := (others => '0');
    variable r4298 : std_logic_vector(0 to 0) := (others => '0');
    variable r4297 : std_logic_vector(0 to 0) := (others => '0');
    variable r4296 : std_logic_vector(0 to 0) := (others => '0');
    variable r4295 : std_logic_vector(0 to 0) := (others => '0');
    variable r4294 : std_logic_vector(0 to 0) := (others => '0');
    variable r4293 : std_logic_vector(0 to 0) := (others => '0');
    variable r4292 : std_logic_vector(0 to 0) := (others => '0');
    variable r4291 : std_logic_vector(0 to 0) := (others => '0');
    variable r4290 : std_logic_vector(0 to 0) := (others => '0');
    variable r4289 : std_logic_vector(0 to 0) := (others => '0');
    variable r4288 : std_logic_vector(0 to 0) := (others => '0');
    variable r4287 : std_logic_vector(0 to 0) := (others => '0');
    variable r4286 : std_logic_vector(0 to 0) := (others => '0');
    variable r4285 : std_logic_vector(0 to 0) := (others => '0');
    variable r4284 : std_logic_vector(0 to 0) := (others => '0');
    variable r4283 : std_logic_vector(0 to 0) := (others => '0');
    variable r4282 : std_logic_vector(0 to 0) := (others => '0');
    variable r4281 : std_logic_vector(0 to 0) := (others => '0');
    variable r4280 : std_logic_vector(0 to 0) := (others => '0');
    variable r4279 : std_logic_vector(0 to 0) := (others => '0');
    variable r4278 : std_logic_vector(0 to 0) := (others => '0');
    variable r4277 : std_logic_vector(0 to 0) := (others => '0');
    variable r4276 : std_logic_vector(0 to 0) := (others => '0');
    variable r4275 : std_logic_vector(0 to 0) := (others => '0');
    variable r4274 : std_logic_vector(0 to 0) := (others => '0');
    variable r4273 : std_logic_vector(0 to 0) := (others => '0');
    variable r4272 : std_logic_vector(0 to 0) := (others => '0');
    variable r4271 : std_logic_vector(0 to 0) := (others => '0');
    variable r4270 : std_logic_vector(0 to 0) := (others => '0');
    variable r4269 : std_logic_vector(0 to 0) := (others => '0');
    variable r4268 : std_logic_vector(0 to 0) := (others => '0');
    variable r4267 : std_logic_vector(0 to 0) := (others => '0');
    variable r4266 : std_logic_vector(0 to 0) := (others => '0');
    variable r4265 : std_logic_vector(0 to 0) := (others => '0');
    variable r4264 : std_logic_vector(0 to 0) := (others => '0');
    variable r4263 : std_logic_vector(0 to 0) := (others => '0');
    variable r4262 : std_logic_vector(0 to 0) := (others => '0');
    variable r4261 : std_logic_vector(0 to 0) := (others => '0');
    variable r4260 : std_logic_vector(0 to 0) := (others => '0');
    variable r4259 : std_logic_vector(0 to 0) := (others => '0');
    variable r4258 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r4259 := "0";
    null;
    r4260 := (r4259);
    r4261 := "0";
    null;
    r4262 := (r4261);
    r4263 := "1";
    null;
    r4264 := (r4263);
    r4265 := "0";
    null;
    r4266 := (r4265);
    r4267 := "1";
    null;
    r4268 := (r4267);
    r4269 := "1";
    null;
    r4270 := (r4269);
    r4271 := "0";
    null;
    r4272 := (r4271);
    r4273 := "1";
    null;
    r4274 := (r4273);
    r4275 := "1";
    null;
    r4276 := (r4275);
    r4277 := "1";
    null;
    r4278 := (r4277);
    r4279 := "1";
    null;
    r4280 := (r4279);
    r4281 := "0";
    null;
    r4282 := (r4281);
    r4283 := "1";
    null;
    r4284 := (r4283);
    r4285 := "0";
    null;
    r4286 := (r4285);
    r4287 := "0";
    null;
    r4288 := (r4287);
    r4289 := "1";
    null;
    r4290 := (r4289);
    r4291 := "0";
    null;
    r4292 := (r4291);
    r4293 := "0";
    null;
    r4294 := (r4293);
    r4295 := "1";
    null;
    r4296 := (r4295);
    r4297 := "0";
    null;
    r4298 := (r4297);
    r4299 := "1";
    null;
    r4300 := (r4299);
    r4301 := "1";
    null;
    r4302 := (r4301);
    r4303 := "0";
    null;
    r4304 := (r4303);
    r4305 := "0";
    null;
    r4306 := (r4305);
    r4307 := "0";
    null;
    r4308 := (r4307);
    r4309 := "1";
    null;
    r4310 := (r4309);
    r4311 := "1";
    null;
    r4312 := (r4311);
    r4313 := "0";
    null;
    r4314 := (r4313);
    r4315 := "1";
    null;
    r4316 := (r4315);
    r4317 := "1";
    null;
    r4318 := (r4317);
    r4319 := "1";
    null;
    r4320 := (r4319);
    r4321 := "1";
    null;
    r4322 := (r4321);
    r4258 := (r4260 & r4262 & r4264 & r4266 & r4268 & r4270 & r4272 & r4274 & r4276 & r4278 & r4280 & r4282 & r4284 & r4286 & r4288 & r4290 & r4292 & r4294 & r4296 & r4298 & r4300 & r4302 & r4304 & r4306 & r4308 & r4310 & r4312 & r4314 & r4316 & r4318 & r4320 & r4322);
    return r4258;
  end rewire_MetaprogrammingRWw2de92c6f_4257;
  function rewire_MetaprogrammingRWw240ca1cc_4188 return std_logic_vector
  is
    variable r4253 : std_logic_vector(0 to 0) := (others => '0');
    variable r4252 : std_logic_vector(0 to 0) := (others => '0');
    variable r4251 : std_logic_vector(0 to 0) := (others => '0');
    variable r4250 : std_logic_vector(0 to 0) := (others => '0');
    variable r4249 : std_logic_vector(0 to 0) := (others => '0');
    variable r4248 : std_logic_vector(0 to 0) := (others => '0');
    variable r4247 : std_logic_vector(0 to 0) := (others => '0');
    variable r4246 : std_logic_vector(0 to 0) := (others => '0');
    variable r4245 : std_logic_vector(0 to 0) := (others => '0');
    variable r4244 : std_logic_vector(0 to 0) := (others => '0');
    variable r4243 : std_logic_vector(0 to 0) := (others => '0');
    variable r4242 : std_logic_vector(0 to 0) := (others => '0');
    variable r4241 : std_logic_vector(0 to 0) := (others => '0');
    variable r4240 : std_logic_vector(0 to 0) := (others => '0');
    variable r4239 : std_logic_vector(0 to 0) := (others => '0');
    variable r4238 : std_logic_vector(0 to 0) := (others => '0');
    variable r4237 : std_logic_vector(0 to 0) := (others => '0');
    variable r4236 : std_logic_vector(0 to 0) := (others => '0');
    variable r4235 : std_logic_vector(0 to 0) := (others => '0');
    variable r4234 : std_logic_vector(0 to 0) := (others => '0');
    variable r4233 : std_logic_vector(0 to 0) := (others => '0');
    variable r4232 : std_logic_vector(0 to 0) := (others => '0');
    variable r4231 : std_logic_vector(0 to 0) := (others => '0');
    variable r4230 : std_logic_vector(0 to 0) := (others => '0');
    variable r4229 : std_logic_vector(0 to 0) := (others => '0');
    variable r4228 : std_logic_vector(0 to 0) := (others => '0');
    variable r4227 : std_logic_vector(0 to 0) := (others => '0');
    variable r4226 : std_logic_vector(0 to 0) := (others => '0');
    variable r4225 : std_logic_vector(0 to 0) := (others => '0');
    variable r4224 : std_logic_vector(0 to 0) := (others => '0');
    variable r4223 : std_logic_vector(0 to 0) := (others => '0');
    variable r4222 : std_logic_vector(0 to 0) := (others => '0');
    variable r4221 : std_logic_vector(0 to 0) := (others => '0');
    variable r4220 : std_logic_vector(0 to 0) := (others => '0');
    variable r4219 : std_logic_vector(0 to 0) := (others => '0');
    variable r4218 : std_logic_vector(0 to 0) := (others => '0');
    variable r4217 : std_logic_vector(0 to 0) := (others => '0');
    variable r4216 : std_logic_vector(0 to 0) := (others => '0');
    variable r4215 : std_logic_vector(0 to 0) := (others => '0');
    variable r4214 : std_logic_vector(0 to 0) := (others => '0');
    variable r4213 : std_logic_vector(0 to 0) := (others => '0');
    variable r4212 : std_logic_vector(0 to 0) := (others => '0');
    variable r4211 : std_logic_vector(0 to 0) := (others => '0');
    variable r4210 : std_logic_vector(0 to 0) := (others => '0');
    variable r4209 : std_logic_vector(0 to 0) := (others => '0');
    variable r4208 : std_logic_vector(0 to 0) := (others => '0');
    variable r4207 : std_logic_vector(0 to 0) := (others => '0');
    variable r4206 : std_logic_vector(0 to 0) := (others => '0');
    variable r4205 : std_logic_vector(0 to 0) := (others => '0');
    variable r4204 : std_logic_vector(0 to 0) := (others => '0');
    variable r4203 : std_logic_vector(0 to 0) := (others => '0');
    variable r4202 : std_logic_vector(0 to 0) := (others => '0');
    variable r4201 : std_logic_vector(0 to 0) := (others => '0');
    variable r4200 : std_logic_vector(0 to 0) := (others => '0');
    variable r4199 : std_logic_vector(0 to 0) := (others => '0');
    variable r4198 : std_logic_vector(0 to 0) := (others => '0');
    variable r4197 : std_logic_vector(0 to 0) := (others => '0');
    variable r4196 : std_logic_vector(0 to 0) := (others => '0');
    variable r4195 : std_logic_vector(0 to 0) := (others => '0');
    variable r4194 : std_logic_vector(0 to 0) := (others => '0');
    variable r4193 : std_logic_vector(0 to 0) := (others => '0');
    variable r4192 : std_logic_vector(0 to 0) := (others => '0');
    variable r4191 : std_logic_vector(0 to 0) := (others => '0');
    variable r4190 : std_logic_vector(0 to 0) := (others => '0');
    variable r4189 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r4190 := "0";
    null;
    r4191 := (r4190);
    r4192 := "0";
    null;
    r4193 := (r4192);
    r4194 := "1";
    null;
    r4195 := (r4194);
    r4196 := "0";
    null;
    r4197 := (r4196);
    r4198 := "0";
    null;
    r4199 := (r4198);
    r4200 := "1";
    null;
    r4201 := (r4200);
    r4202 := "0";
    null;
    r4203 := (r4202);
    r4204 := "0";
    null;
    r4205 := (r4204);
    r4206 := "0";
    null;
    r4207 := (r4206);
    r4208 := "0";
    null;
    r4209 := (r4208);
    r4210 := "0";
    null;
    r4211 := (r4210);
    r4212 := "0";
    null;
    r4213 := (r4212);
    r4214 := "1";
    null;
    r4215 := (r4214);
    r4216 := "1";
    null;
    r4217 := (r4216);
    r4218 := "0";
    null;
    r4219 := (r4218);
    r4220 := "0";
    null;
    r4221 := (r4220);
    r4222 := "1";
    null;
    r4223 := (r4222);
    r4224 := "0";
    null;
    r4225 := (r4224);
    r4226 := "1";
    null;
    r4227 := (r4226);
    r4228 := "0";
    null;
    r4229 := (r4228);
    r4230 := "0";
    null;
    r4231 := (r4230);
    r4232 := "0";
    null;
    r4233 := (r4232);
    r4234 := "0";
    null;
    r4235 := (r4234);
    r4236 := "1";
    null;
    r4237 := (r4236);
    r4238 := "1";
    null;
    r4239 := (r4238);
    r4240 := "1";
    null;
    r4241 := (r4240);
    r4242 := "0";
    null;
    r4243 := (r4242);
    r4244 := "0";
    null;
    r4245 := (r4244);
    r4246 := "1";
    null;
    r4247 := (r4246);
    r4248 := "1";
    null;
    r4249 := (r4248);
    r4250 := "0";
    null;
    r4251 := (r4250);
    r4252 := "0";
    null;
    r4253 := (r4252);
    r4189 := (r4191 & r4193 & r4195 & r4197 & r4199 & r4201 & r4203 & r4205 & r4207 & r4209 & r4211 & r4213 & r4215 & r4217 & r4219 & r4221 & r4223 & r4225 & r4227 & r4229 & r4231 & r4233 & r4235 & r4237 & r4239 & r4241 & r4243 & r4245 & r4247 & r4249 & r4251 & r4253);
    return r4189;
  end rewire_MetaprogrammingRWw240ca1cc_4188;
  function rewire_MetaprogrammingRWw0fc19dc6_4119 return std_logic_vector
  is
    variable r4184 : std_logic_vector(0 to 0) := (others => '0');
    variable r4183 : std_logic_vector(0 to 0) := (others => '0');
    variable r4182 : std_logic_vector(0 to 0) := (others => '0');
    variable r4181 : std_logic_vector(0 to 0) := (others => '0');
    variable r4180 : std_logic_vector(0 to 0) := (others => '0');
    variable r4179 : std_logic_vector(0 to 0) := (others => '0');
    variable r4178 : std_logic_vector(0 to 0) := (others => '0');
    variable r4177 : std_logic_vector(0 to 0) := (others => '0');
    variable r4176 : std_logic_vector(0 to 0) := (others => '0');
    variable r4175 : std_logic_vector(0 to 0) := (others => '0');
    variable r4174 : std_logic_vector(0 to 0) := (others => '0');
    variable r4173 : std_logic_vector(0 to 0) := (others => '0');
    variable r4172 : std_logic_vector(0 to 0) := (others => '0');
    variable r4171 : std_logic_vector(0 to 0) := (others => '0');
    variable r4170 : std_logic_vector(0 to 0) := (others => '0');
    variable r4169 : std_logic_vector(0 to 0) := (others => '0');
    variable r4168 : std_logic_vector(0 to 0) := (others => '0');
    variable r4167 : std_logic_vector(0 to 0) := (others => '0');
    variable r4166 : std_logic_vector(0 to 0) := (others => '0');
    variable r4165 : std_logic_vector(0 to 0) := (others => '0');
    variable r4164 : std_logic_vector(0 to 0) := (others => '0');
    variable r4163 : std_logic_vector(0 to 0) := (others => '0');
    variable r4162 : std_logic_vector(0 to 0) := (others => '0');
    variable r4161 : std_logic_vector(0 to 0) := (others => '0');
    variable r4160 : std_logic_vector(0 to 0) := (others => '0');
    variable r4159 : std_logic_vector(0 to 0) := (others => '0');
    variable r4158 : std_logic_vector(0 to 0) := (others => '0');
    variable r4157 : std_logic_vector(0 to 0) := (others => '0');
    variable r4156 : std_logic_vector(0 to 0) := (others => '0');
    variable r4155 : std_logic_vector(0 to 0) := (others => '0');
    variable r4154 : std_logic_vector(0 to 0) := (others => '0');
    variable r4153 : std_logic_vector(0 to 0) := (others => '0');
    variable r4152 : std_logic_vector(0 to 0) := (others => '0');
    variable r4151 : std_logic_vector(0 to 0) := (others => '0');
    variable r4150 : std_logic_vector(0 to 0) := (others => '0');
    variable r4149 : std_logic_vector(0 to 0) := (others => '0');
    variable r4148 : std_logic_vector(0 to 0) := (others => '0');
    variable r4147 : std_logic_vector(0 to 0) := (others => '0');
    variable r4146 : std_logic_vector(0 to 0) := (others => '0');
    variable r4145 : std_logic_vector(0 to 0) := (others => '0');
    variable r4144 : std_logic_vector(0 to 0) := (others => '0');
    variable r4143 : std_logic_vector(0 to 0) := (others => '0');
    variable r4142 : std_logic_vector(0 to 0) := (others => '0');
    variable r4141 : std_logic_vector(0 to 0) := (others => '0');
    variable r4140 : std_logic_vector(0 to 0) := (others => '0');
    variable r4139 : std_logic_vector(0 to 0) := (others => '0');
    variable r4138 : std_logic_vector(0 to 0) := (others => '0');
    variable r4137 : std_logic_vector(0 to 0) := (others => '0');
    variable r4136 : std_logic_vector(0 to 0) := (others => '0');
    variable r4135 : std_logic_vector(0 to 0) := (others => '0');
    variable r4134 : std_logic_vector(0 to 0) := (others => '0');
    variable r4133 : std_logic_vector(0 to 0) := (others => '0');
    variable r4132 : std_logic_vector(0 to 0) := (others => '0');
    variable r4131 : std_logic_vector(0 to 0) := (others => '0');
    variable r4130 : std_logic_vector(0 to 0) := (others => '0');
    variable r4129 : std_logic_vector(0 to 0) := (others => '0');
    variable r4128 : std_logic_vector(0 to 0) := (others => '0');
    variable r4127 : std_logic_vector(0 to 0) := (others => '0');
    variable r4126 : std_logic_vector(0 to 0) := (others => '0');
    variable r4125 : std_logic_vector(0 to 0) := (others => '0');
    variable r4124 : std_logic_vector(0 to 0) := (others => '0');
    variable r4123 : std_logic_vector(0 to 0) := (others => '0');
    variable r4122 : std_logic_vector(0 to 0) := (others => '0');
    variable r4121 : std_logic_vector(0 to 0) := (others => '0');
    variable r4120 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r4121 := "0";
    null;
    r4122 := (r4121);
    r4123 := "0";
    null;
    r4124 := (r4123);
    r4125 := "0";
    null;
    r4126 := (r4125);
    r4127 := "0";
    null;
    r4128 := (r4127);
    r4129 := "1";
    null;
    r4130 := (r4129);
    r4131 := "1";
    null;
    r4132 := (r4131);
    r4133 := "1";
    null;
    r4134 := (r4133);
    r4135 := "1";
    null;
    r4136 := (r4135);
    r4137 := "1";
    null;
    r4138 := (r4137);
    r4139 := "1";
    null;
    r4140 := (r4139);
    r4141 := "0";
    null;
    r4142 := (r4141);
    r4143 := "0";
    null;
    r4144 := (r4143);
    r4145 := "0";
    null;
    r4146 := (r4145);
    r4147 := "0";
    null;
    r4148 := (r4147);
    r4149 := "0";
    null;
    r4150 := (r4149);
    r4151 := "1";
    null;
    r4152 := (r4151);
    r4153 := "1";
    null;
    r4154 := (r4153);
    r4155 := "0";
    null;
    r4156 := (r4155);
    r4157 := "0";
    null;
    r4158 := (r4157);
    r4159 := "1";
    null;
    r4160 := (r4159);
    r4161 := "1";
    null;
    r4162 := (r4161);
    r4163 := "1";
    null;
    r4164 := (r4163);
    r4165 := "0";
    null;
    r4166 := (r4165);
    r4167 := "1";
    null;
    r4168 := (r4167);
    r4169 := "1";
    null;
    r4170 := (r4169);
    r4171 := "1";
    null;
    r4172 := (r4171);
    r4173 := "0";
    null;
    r4174 := (r4173);
    r4175 := "0";
    null;
    r4176 := (r4175);
    r4177 := "0";
    null;
    r4178 := (r4177);
    r4179 := "1";
    null;
    r4180 := (r4179);
    r4181 := "1";
    null;
    r4182 := (r4181);
    r4183 := "0";
    null;
    r4184 := (r4183);
    r4120 := (r4122 & r4124 & r4126 & r4128 & r4130 & r4132 & r4134 & r4136 & r4138 & r4140 & r4142 & r4144 & r4146 & r4148 & r4150 & r4152 & r4154 & r4156 & r4158 & r4160 & r4162 & r4164 & r4166 & r4168 & r4170 & r4172 & r4174 & r4176 & r4178 & r4180 & r4182 & r4184);
    return r4120;
  end rewire_MetaprogrammingRWw0fc19dc6_4119;
  function rewire_MetaprogrammingRWwefbe4786_4050 return std_logic_vector
  is
    variable r4115 : std_logic_vector(0 to 0) := (others => '0');
    variable r4114 : std_logic_vector(0 to 0) := (others => '0');
    variable r4113 : std_logic_vector(0 to 0) := (others => '0');
    variable r4112 : std_logic_vector(0 to 0) := (others => '0');
    variable r4111 : std_logic_vector(0 to 0) := (others => '0');
    variable r4110 : std_logic_vector(0 to 0) := (others => '0');
    variable r4109 : std_logic_vector(0 to 0) := (others => '0');
    variable r4108 : std_logic_vector(0 to 0) := (others => '0');
    variable r4107 : std_logic_vector(0 to 0) := (others => '0');
    variable r4106 : std_logic_vector(0 to 0) := (others => '0');
    variable r4105 : std_logic_vector(0 to 0) := (others => '0');
    variable r4104 : std_logic_vector(0 to 0) := (others => '0');
    variable r4103 : std_logic_vector(0 to 0) := (others => '0');
    variable r4102 : std_logic_vector(0 to 0) := (others => '0');
    variable r4101 : std_logic_vector(0 to 0) := (others => '0');
    variable r4100 : std_logic_vector(0 to 0) := (others => '0');
    variable r4099 : std_logic_vector(0 to 0) := (others => '0');
    variable r4098 : std_logic_vector(0 to 0) := (others => '0');
    variable r4097 : std_logic_vector(0 to 0) := (others => '0');
    variable r4096 : std_logic_vector(0 to 0) := (others => '0');
    variable r4095 : std_logic_vector(0 to 0) := (others => '0');
    variable r4094 : std_logic_vector(0 to 0) := (others => '0');
    variable r4093 : std_logic_vector(0 to 0) := (others => '0');
    variable r4092 : std_logic_vector(0 to 0) := (others => '0');
    variable r4091 : std_logic_vector(0 to 0) := (others => '0');
    variable r4090 : std_logic_vector(0 to 0) := (others => '0');
    variable r4089 : std_logic_vector(0 to 0) := (others => '0');
    variable r4088 : std_logic_vector(0 to 0) := (others => '0');
    variable r4087 : std_logic_vector(0 to 0) := (others => '0');
    variable r4086 : std_logic_vector(0 to 0) := (others => '0');
    variable r4085 : std_logic_vector(0 to 0) := (others => '0');
    variable r4084 : std_logic_vector(0 to 0) := (others => '0');
    variable r4083 : std_logic_vector(0 to 0) := (others => '0');
    variable r4082 : std_logic_vector(0 to 0) := (others => '0');
    variable r4081 : std_logic_vector(0 to 0) := (others => '0');
    variable r4080 : std_logic_vector(0 to 0) := (others => '0');
    variable r4079 : std_logic_vector(0 to 0) := (others => '0');
    variable r4078 : std_logic_vector(0 to 0) := (others => '0');
    variable r4077 : std_logic_vector(0 to 0) := (others => '0');
    variable r4076 : std_logic_vector(0 to 0) := (others => '0');
    variable r4075 : std_logic_vector(0 to 0) := (others => '0');
    variable r4074 : std_logic_vector(0 to 0) := (others => '0');
    variable r4073 : std_logic_vector(0 to 0) := (others => '0');
    variable r4072 : std_logic_vector(0 to 0) := (others => '0');
    variable r4071 : std_logic_vector(0 to 0) := (others => '0');
    variable r4070 : std_logic_vector(0 to 0) := (others => '0');
    variable r4069 : std_logic_vector(0 to 0) := (others => '0');
    variable r4068 : std_logic_vector(0 to 0) := (others => '0');
    variable r4067 : std_logic_vector(0 to 0) := (others => '0');
    variable r4066 : std_logic_vector(0 to 0) := (others => '0');
    variable r4065 : std_logic_vector(0 to 0) := (others => '0');
    variable r4064 : std_logic_vector(0 to 0) := (others => '0');
    variable r4063 : std_logic_vector(0 to 0) := (others => '0');
    variable r4062 : std_logic_vector(0 to 0) := (others => '0');
    variable r4061 : std_logic_vector(0 to 0) := (others => '0');
    variable r4060 : std_logic_vector(0 to 0) := (others => '0');
    variable r4059 : std_logic_vector(0 to 0) := (others => '0');
    variable r4058 : std_logic_vector(0 to 0) := (others => '0');
    variable r4057 : std_logic_vector(0 to 0) := (others => '0');
    variable r4056 : std_logic_vector(0 to 0) := (others => '0');
    variable r4055 : std_logic_vector(0 to 0) := (others => '0');
    variable r4054 : std_logic_vector(0 to 0) := (others => '0');
    variable r4053 : std_logic_vector(0 to 0) := (others => '0');
    variable r4052 : std_logic_vector(0 to 0) := (others => '0');
    variable r4051 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r4052 := "1";
    null;
    r4053 := (r4052);
    r4054 := "1";
    null;
    r4055 := (r4054);
    r4056 := "1";
    null;
    r4057 := (r4056);
    r4058 := "0";
    null;
    r4059 := (r4058);
    r4060 := "1";
    null;
    r4061 := (r4060);
    r4062 := "1";
    null;
    r4063 := (r4062);
    r4064 := "1";
    null;
    r4065 := (r4064);
    r4066 := "1";
    null;
    r4067 := (r4066);
    r4068 := "1";
    null;
    r4069 := (r4068);
    r4070 := "0";
    null;
    r4071 := (r4070);
    r4072 := "1";
    null;
    r4073 := (r4072);
    r4074 := "1";
    null;
    r4075 := (r4074);
    r4076 := "1";
    null;
    r4077 := (r4076);
    r4078 := "1";
    null;
    r4079 := (r4078);
    r4080 := "1";
    null;
    r4081 := (r4080);
    r4082 := "0";
    null;
    r4083 := (r4082);
    r4084 := "0";
    null;
    r4085 := (r4084);
    r4086 := "1";
    null;
    r4087 := (r4086);
    r4088 := "0";
    null;
    r4089 := (r4088);
    r4090 := "0";
    null;
    r4091 := (r4090);
    r4092 := "0";
    null;
    r4093 := (r4092);
    r4094 := "1";
    null;
    r4095 := (r4094);
    r4096 := "1";
    null;
    r4097 := (r4096);
    r4098 := "1";
    null;
    r4099 := (r4098);
    r4100 := "1";
    null;
    r4101 := (r4100);
    r4102 := "0";
    null;
    r4103 := (r4102);
    r4104 := "0";
    null;
    r4105 := (r4104);
    r4106 := "0";
    null;
    r4107 := (r4106);
    r4108 := "0";
    null;
    r4109 := (r4108);
    r4110 := "1";
    null;
    r4111 := (r4110);
    r4112 := "1";
    null;
    r4113 := (r4112);
    r4114 := "0";
    null;
    r4115 := (r4114);
    r4051 := (r4053 & r4055 & r4057 & r4059 & r4061 & r4063 & r4065 & r4067 & r4069 & r4071 & r4073 & r4075 & r4077 & r4079 & r4081 & r4083 & r4085 & r4087 & r4089 & r4091 & r4093 & r4095 & r4097 & r4099 & r4101 & r4103 & r4105 & r4107 & r4109 & r4111 & r4113 & r4115);
    return r4051;
  end rewire_MetaprogrammingRWwefbe4786_4050;
  function rewire_MetaprogrammingRWwe49b69c1_3981 return std_logic_vector
  is
    variable r4046 : std_logic_vector(0 to 0) := (others => '0');
    variable r4045 : std_logic_vector(0 to 0) := (others => '0');
    variable r4044 : std_logic_vector(0 to 0) := (others => '0');
    variable r4043 : std_logic_vector(0 to 0) := (others => '0');
    variable r4042 : std_logic_vector(0 to 0) := (others => '0');
    variable r4041 : std_logic_vector(0 to 0) := (others => '0');
    variable r4040 : std_logic_vector(0 to 0) := (others => '0');
    variable r4039 : std_logic_vector(0 to 0) := (others => '0');
    variable r4038 : std_logic_vector(0 to 0) := (others => '0');
    variable r4037 : std_logic_vector(0 to 0) := (others => '0');
    variable r4036 : std_logic_vector(0 to 0) := (others => '0');
    variable r4035 : std_logic_vector(0 to 0) := (others => '0');
    variable r4034 : std_logic_vector(0 to 0) := (others => '0');
    variable r4033 : std_logic_vector(0 to 0) := (others => '0');
    variable r4032 : std_logic_vector(0 to 0) := (others => '0');
    variable r4031 : std_logic_vector(0 to 0) := (others => '0');
    variable r4030 : std_logic_vector(0 to 0) := (others => '0');
    variable r4029 : std_logic_vector(0 to 0) := (others => '0');
    variable r4028 : std_logic_vector(0 to 0) := (others => '0');
    variable r4027 : std_logic_vector(0 to 0) := (others => '0');
    variable r4026 : std_logic_vector(0 to 0) := (others => '0');
    variable r4025 : std_logic_vector(0 to 0) := (others => '0');
    variable r4024 : std_logic_vector(0 to 0) := (others => '0');
    variable r4023 : std_logic_vector(0 to 0) := (others => '0');
    variable r4022 : std_logic_vector(0 to 0) := (others => '0');
    variable r4021 : std_logic_vector(0 to 0) := (others => '0');
    variable r4020 : std_logic_vector(0 to 0) := (others => '0');
    variable r4019 : std_logic_vector(0 to 0) := (others => '0');
    variable r4018 : std_logic_vector(0 to 0) := (others => '0');
    variable r4017 : std_logic_vector(0 to 0) := (others => '0');
    variable r4016 : std_logic_vector(0 to 0) := (others => '0');
    variable r4015 : std_logic_vector(0 to 0) := (others => '0');
    variable r4014 : std_logic_vector(0 to 0) := (others => '0');
    variable r4013 : std_logic_vector(0 to 0) := (others => '0');
    variable r4012 : std_logic_vector(0 to 0) := (others => '0');
    variable r4011 : std_logic_vector(0 to 0) := (others => '0');
    variable r4010 : std_logic_vector(0 to 0) := (others => '0');
    variable r4009 : std_logic_vector(0 to 0) := (others => '0');
    variable r4008 : std_logic_vector(0 to 0) := (others => '0');
    variable r4007 : std_logic_vector(0 to 0) := (others => '0');
    variable r4006 : std_logic_vector(0 to 0) := (others => '0');
    variable r4005 : std_logic_vector(0 to 0) := (others => '0');
    variable r4004 : std_logic_vector(0 to 0) := (others => '0');
    variable r4003 : std_logic_vector(0 to 0) := (others => '0');
    variable r4002 : std_logic_vector(0 to 0) := (others => '0');
    variable r4001 : std_logic_vector(0 to 0) := (others => '0');
    variable r4000 : std_logic_vector(0 to 0) := (others => '0');
    variable r3999 : std_logic_vector(0 to 0) := (others => '0');
    variable r3998 : std_logic_vector(0 to 0) := (others => '0');
    variable r3997 : std_logic_vector(0 to 0) := (others => '0');
    variable r3996 : std_logic_vector(0 to 0) := (others => '0');
    variable r3995 : std_logic_vector(0 to 0) := (others => '0');
    variable r3994 : std_logic_vector(0 to 0) := (others => '0');
    variable r3993 : std_logic_vector(0 to 0) := (others => '0');
    variable r3992 : std_logic_vector(0 to 0) := (others => '0');
    variable r3991 : std_logic_vector(0 to 0) := (others => '0');
    variable r3990 : std_logic_vector(0 to 0) := (others => '0');
    variable r3989 : std_logic_vector(0 to 0) := (others => '0');
    variable r3988 : std_logic_vector(0 to 0) := (others => '0');
    variable r3987 : std_logic_vector(0 to 0) := (others => '0');
    variable r3986 : std_logic_vector(0 to 0) := (others => '0');
    variable r3985 : std_logic_vector(0 to 0) := (others => '0');
    variable r3984 : std_logic_vector(0 to 0) := (others => '0');
    variable r3983 : std_logic_vector(0 to 0) := (others => '0');
    variable r3982 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r3983 := "1";
    null;
    r3984 := (r3983);
    r3985 := "1";
    null;
    r3986 := (r3985);
    r3987 := "1";
    null;
    r3988 := (r3987);
    r3989 := "0";
    null;
    r3990 := (r3989);
    r3991 := "0";
    null;
    r3992 := (r3991);
    r3993 := "1";
    null;
    r3994 := (r3993);
    r3995 := "0";
    null;
    r3996 := (r3995);
    r3997 := "0";
    null;
    r3998 := (r3997);
    r3999 := "1";
    null;
    r4000 := (r3999);
    r4001 := "0";
    null;
    r4002 := (r4001);
    r4003 := "0";
    null;
    r4004 := (r4003);
    r4005 := "1";
    null;
    r4006 := (r4005);
    r4007 := "1";
    null;
    r4008 := (r4007);
    r4009 := "0";
    null;
    r4010 := (r4009);
    r4011 := "1";
    null;
    r4012 := (r4011);
    r4013 := "1";
    null;
    r4014 := (r4013);
    r4015 := "0";
    null;
    r4016 := (r4015);
    r4017 := "1";
    null;
    r4018 := (r4017);
    r4019 := "1";
    null;
    r4020 := (r4019);
    r4021 := "0";
    null;
    r4022 := (r4021);
    r4023 := "1";
    null;
    r4024 := (r4023);
    r4025 := "0";
    null;
    r4026 := (r4025);
    r4027 := "0";
    null;
    r4028 := (r4027);
    r4029 := "1";
    null;
    r4030 := (r4029);
    r4031 := "1";
    null;
    r4032 := (r4031);
    r4033 := "1";
    null;
    r4034 := (r4033);
    r4035 := "0";
    null;
    r4036 := (r4035);
    r4037 := "0";
    null;
    r4038 := (r4037);
    r4039 := "0";
    null;
    r4040 := (r4039);
    r4041 := "0";
    null;
    r4042 := (r4041);
    r4043 := "0";
    null;
    r4044 := (r4043);
    r4045 := "1";
    null;
    r4046 := (r4045);
    r3982 := (r3984 & r3986 & r3988 & r3990 & r3992 & r3994 & r3996 & r3998 & r4000 & r4002 & r4004 & r4006 & r4008 & r4010 & r4012 & r4014 & r4016 & r4018 & r4020 & r4022 & r4024 & r4026 & r4028 & r4030 & r4032 & r4034 & r4036 & r4038 & r4040 & r4042 & r4044 & r4046);
    return r3982;
  end rewire_MetaprogrammingRWwe49b69c1_3981;
  function rewire_MetaprogrammingRWwc19bf174_3912 return std_logic_vector
  is
    variable r3977 : std_logic_vector(0 to 0) := (others => '0');
    variable r3976 : std_logic_vector(0 to 0) := (others => '0');
    variable r3975 : std_logic_vector(0 to 0) := (others => '0');
    variable r3974 : std_logic_vector(0 to 0) := (others => '0');
    variable r3973 : std_logic_vector(0 to 0) := (others => '0');
    variable r3972 : std_logic_vector(0 to 0) := (others => '0');
    variable r3971 : std_logic_vector(0 to 0) := (others => '0');
    variable r3970 : std_logic_vector(0 to 0) := (others => '0');
    variable r3969 : std_logic_vector(0 to 0) := (others => '0');
    variable r3968 : std_logic_vector(0 to 0) := (others => '0');
    variable r3967 : std_logic_vector(0 to 0) := (others => '0');
    variable r3966 : std_logic_vector(0 to 0) := (others => '0');
    variable r3965 : std_logic_vector(0 to 0) := (others => '0');
    variable r3964 : std_logic_vector(0 to 0) := (others => '0');
    variable r3963 : std_logic_vector(0 to 0) := (others => '0');
    variable r3962 : std_logic_vector(0 to 0) := (others => '0');
    variable r3961 : std_logic_vector(0 to 0) := (others => '0');
    variable r3960 : std_logic_vector(0 to 0) := (others => '0');
    variable r3959 : std_logic_vector(0 to 0) := (others => '0');
    variable r3958 : std_logic_vector(0 to 0) := (others => '0');
    variable r3957 : std_logic_vector(0 to 0) := (others => '0');
    variable r3956 : std_logic_vector(0 to 0) := (others => '0');
    variable r3955 : std_logic_vector(0 to 0) := (others => '0');
    variable r3954 : std_logic_vector(0 to 0) := (others => '0');
    variable r3953 : std_logic_vector(0 to 0) := (others => '0');
    variable r3952 : std_logic_vector(0 to 0) := (others => '0');
    variable r3951 : std_logic_vector(0 to 0) := (others => '0');
    variable r3950 : std_logic_vector(0 to 0) := (others => '0');
    variable r3949 : std_logic_vector(0 to 0) := (others => '0');
    variable r3948 : std_logic_vector(0 to 0) := (others => '0');
    variable r3947 : std_logic_vector(0 to 0) := (others => '0');
    variable r3946 : std_logic_vector(0 to 0) := (others => '0');
    variable r3945 : std_logic_vector(0 to 0) := (others => '0');
    variable r3944 : std_logic_vector(0 to 0) := (others => '0');
    variable r3943 : std_logic_vector(0 to 0) := (others => '0');
    variable r3942 : std_logic_vector(0 to 0) := (others => '0');
    variable r3941 : std_logic_vector(0 to 0) := (others => '0');
    variable r3940 : std_logic_vector(0 to 0) := (others => '0');
    variable r3939 : std_logic_vector(0 to 0) := (others => '0');
    variable r3938 : std_logic_vector(0 to 0) := (others => '0');
    variable r3937 : std_logic_vector(0 to 0) := (others => '0');
    variable r3936 : std_logic_vector(0 to 0) := (others => '0');
    variable r3935 : std_logic_vector(0 to 0) := (others => '0');
    variable r3934 : std_logic_vector(0 to 0) := (others => '0');
    variable r3933 : std_logic_vector(0 to 0) := (others => '0');
    variable r3932 : std_logic_vector(0 to 0) := (others => '0');
    variable r3931 : std_logic_vector(0 to 0) := (others => '0');
    variable r3930 : std_logic_vector(0 to 0) := (others => '0');
    variable r3929 : std_logic_vector(0 to 0) := (others => '0');
    variable r3928 : std_logic_vector(0 to 0) := (others => '0');
    variable r3927 : std_logic_vector(0 to 0) := (others => '0');
    variable r3926 : std_logic_vector(0 to 0) := (others => '0');
    variable r3925 : std_logic_vector(0 to 0) := (others => '0');
    variable r3924 : std_logic_vector(0 to 0) := (others => '0');
    variable r3923 : std_logic_vector(0 to 0) := (others => '0');
    variable r3922 : std_logic_vector(0 to 0) := (others => '0');
    variable r3921 : std_logic_vector(0 to 0) := (others => '0');
    variable r3920 : std_logic_vector(0 to 0) := (others => '0');
    variable r3919 : std_logic_vector(0 to 0) := (others => '0');
    variable r3918 : std_logic_vector(0 to 0) := (others => '0');
    variable r3917 : std_logic_vector(0 to 0) := (others => '0');
    variable r3916 : std_logic_vector(0 to 0) := (others => '0');
    variable r3915 : std_logic_vector(0 to 0) := (others => '0');
    variable r3914 : std_logic_vector(0 to 0) := (others => '0');
    variable r3913 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r3914 := "1";
    null;
    r3915 := (r3914);
    r3916 := "1";
    null;
    r3917 := (r3916);
    r3918 := "0";
    null;
    r3919 := (r3918);
    r3920 := "0";
    null;
    r3921 := (r3920);
    r3922 := "0";
    null;
    r3923 := (r3922);
    r3924 := "0";
    null;
    r3925 := (r3924);
    r3926 := "0";
    null;
    r3927 := (r3926);
    r3928 := "1";
    null;
    r3929 := (r3928);
    r3930 := "1";
    null;
    r3931 := (r3930);
    r3932 := "0";
    null;
    r3933 := (r3932);
    r3934 := "0";
    null;
    r3935 := (r3934);
    r3936 := "1";
    null;
    r3937 := (r3936);
    r3938 := "1";
    null;
    r3939 := (r3938);
    r3940 := "0";
    null;
    r3941 := (r3940);
    r3942 := "1";
    null;
    r3943 := (r3942);
    r3944 := "1";
    null;
    r3945 := (r3944);
    r3946 := "1";
    null;
    r3947 := (r3946);
    r3948 := "1";
    null;
    r3949 := (r3948);
    r3950 := "1";
    null;
    r3951 := (r3950);
    r3952 := "1";
    null;
    r3953 := (r3952);
    r3954 := "0";
    null;
    r3955 := (r3954);
    r3956 := "0";
    null;
    r3957 := (r3956);
    r3958 := "0";
    null;
    r3959 := (r3958);
    r3960 := "1";
    null;
    r3961 := (r3960);
    r3962 := "0";
    null;
    r3963 := (r3962);
    r3964 := "1";
    null;
    r3965 := (r3964);
    r3966 := "1";
    null;
    r3967 := (r3966);
    r3968 := "1";
    null;
    r3969 := (r3968);
    r3970 := "0";
    null;
    r3971 := (r3970);
    r3972 := "1";
    null;
    r3973 := (r3972);
    r3974 := "0";
    null;
    r3975 := (r3974);
    r3976 := "0";
    null;
    r3977 := (r3976);
    r3913 := (r3915 & r3917 & r3919 & r3921 & r3923 & r3925 & r3927 & r3929 & r3931 & r3933 & r3935 & r3937 & r3939 & r3941 & r3943 & r3945 & r3947 & r3949 & r3951 & r3953 & r3955 & r3957 & r3959 & r3961 & r3963 & r3965 & r3967 & r3969 & r3971 & r3973 & r3975 & r3977);
    return r3913;
  end rewire_MetaprogrammingRWwc19bf174_3912;
  function rewire_MetaprogrammingRWw9bdc06a7_3843 return std_logic_vector
  is
    variable r3908 : std_logic_vector(0 to 0) := (others => '0');
    variable r3907 : std_logic_vector(0 to 0) := (others => '0');
    variable r3906 : std_logic_vector(0 to 0) := (others => '0');
    variable r3905 : std_logic_vector(0 to 0) := (others => '0');
    variable r3904 : std_logic_vector(0 to 0) := (others => '0');
    variable r3903 : std_logic_vector(0 to 0) := (others => '0');
    variable r3902 : std_logic_vector(0 to 0) := (others => '0');
    variable r3901 : std_logic_vector(0 to 0) := (others => '0');
    variable r3900 : std_logic_vector(0 to 0) := (others => '0');
    variable r3899 : std_logic_vector(0 to 0) := (others => '0');
    variable r3898 : std_logic_vector(0 to 0) := (others => '0');
    variable r3897 : std_logic_vector(0 to 0) := (others => '0');
    variable r3896 : std_logic_vector(0 to 0) := (others => '0');
    variable r3895 : std_logic_vector(0 to 0) := (others => '0');
    variable r3894 : std_logic_vector(0 to 0) := (others => '0');
    variable r3893 : std_logic_vector(0 to 0) := (others => '0');
    variable r3892 : std_logic_vector(0 to 0) := (others => '0');
    variable r3891 : std_logic_vector(0 to 0) := (others => '0');
    variable r3890 : std_logic_vector(0 to 0) := (others => '0');
    variable r3889 : std_logic_vector(0 to 0) := (others => '0');
    variable r3888 : std_logic_vector(0 to 0) := (others => '0');
    variable r3887 : std_logic_vector(0 to 0) := (others => '0');
    variable r3886 : std_logic_vector(0 to 0) := (others => '0');
    variable r3885 : std_logic_vector(0 to 0) := (others => '0');
    variable r3884 : std_logic_vector(0 to 0) := (others => '0');
    variable r3883 : std_logic_vector(0 to 0) := (others => '0');
    variable r3882 : std_logic_vector(0 to 0) := (others => '0');
    variable r3881 : std_logic_vector(0 to 0) := (others => '0');
    variable r3880 : std_logic_vector(0 to 0) := (others => '0');
    variable r3879 : std_logic_vector(0 to 0) := (others => '0');
    variable r3878 : std_logic_vector(0 to 0) := (others => '0');
    variable r3877 : std_logic_vector(0 to 0) := (others => '0');
    variable r3876 : std_logic_vector(0 to 0) := (others => '0');
    variable r3875 : std_logic_vector(0 to 0) := (others => '0');
    variable r3874 : std_logic_vector(0 to 0) := (others => '0');
    variable r3873 : std_logic_vector(0 to 0) := (others => '0');
    variable r3872 : std_logic_vector(0 to 0) := (others => '0');
    variable r3871 : std_logic_vector(0 to 0) := (others => '0');
    variable r3870 : std_logic_vector(0 to 0) := (others => '0');
    variable r3869 : std_logic_vector(0 to 0) := (others => '0');
    variable r3868 : std_logic_vector(0 to 0) := (others => '0');
    variable r3867 : std_logic_vector(0 to 0) := (others => '0');
    variable r3866 : std_logic_vector(0 to 0) := (others => '0');
    variable r3865 : std_logic_vector(0 to 0) := (others => '0');
    variable r3864 : std_logic_vector(0 to 0) := (others => '0');
    variable r3863 : std_logic_vector(0 to 0) := (others => '0');
    variable r3862 : std_logic_vector(0 to 0) := (others => '0');
    variable r3861 : std_logic_vector(0 to 0) := (others => '0');
    variable r3860 : std_logic_vector(0 to 0) := (others => '0');
    variable r3859 : std_logic_vector(0 to 0) := (others => '0');
    variable r3858 : std_logic_vector(0 to 0) := (others => '0');
    variable r3857 : std_logic_vector(0 to 0) := (others => '0');
    variable r3856 : std_logic_vector(0 to 0) := (others => '0');
    variable r3855 : std_logic_vector(0 to 0) := (others => '0');
    variable r3854 : std_logic_vector(0 to 0) := (others => '0');
    variable r3853 : std_logic_vector(0 to 0) := (others => '0');
    variable r3852 : std_logic_vector(0 to 0) := (others => '0');
    variable r3851 : std_logic_vector(0 to 0) := (others => '0');
    variable r3850 : std_logic_vector(0 to 0) := (others => '0');
    variable r3849 : std_logic_vector(0 to 0) := (others => '0');
    variable r3848 : std_logic_vector(0 to 0) := (others => '0');
    variable r3847 : std_logic_vector(0 to 0) := (others => '0');
    variable r3846 : std_logic_vector(0 to 0) := (others => '0');
    variable r3845 : std_logic_vector(0 to 0) := (others => '0');
    variable r3844 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r3845 := "1";
    null;
    r3846 := (r3845);
    r3847 := "0";
    null;
    r3848 := (r3847);
    r3849 := "0";
    null;
    r3850 := (r3849);
    r3851 := "1";
    null;
    r3852 := (r3851);
    r3853 := "1";
    null;
    r3854 := (r3853);
    r3855 := "0";
    null;
    r3856 := (r3855);
    r3857 := "1";
    null;
    r3858 := (r3857);
    r3859 := "1";
    null;
    r3860 := (r3859);
    r3861 := "1";
    null;
    r3862 := (r3861);
    r3863 := "1";
    null;
    r3864 := (r3863);
    r3865 := "0";
    null;
    r3866 := (r3865);
    r3867 := "1";
    null;
    r3868 := (r3867);
    r3869 := "1";
    null;
    r3870 := (r3869);
    r3871 := "1";
    null;
    r3872 := (r3871);
    r3873 := "0";
    null;
    r3874 := (r3873);
    r3875 := "0";
    null;
    r3876 := (r3875);
    r3877 := "0";
    null;
    r3878 := (r3877);
    r3879 := "0";
    null;
    r3880 := (r3879);
    r3881 := "0";
    null;
    r3882 := (r3881);
    r3883 := "0";
    null;
    r3884 := (r3883);
    r3885 := "0";
    null;
    r3886 := (r3885);
    r3887 := "1";
    null;
    r3888 := (r3887);
    r3889 := "1";
    null;
    r3890 := (r3889);
    r3891 := "0";
    null;
    r3892 := (r3891);
    r3893 := "1";
    null;
    r3894 := (r3893);
    r3895 := "0";
    null;
    r3896 := (r3895);
    r3897 := "1";
    null;
    r3898 := (r3897);
    r3899 := "0";
    null;
    r3900 := (r3899);
    r3901 := "0";
    null;
    r3902 := (r3901);
    r3903 := "1";
    null;
    r3904 := (r3903);
    r3905 := "1";
    null;
    r3906 := (r3905);
    r3907 := "1";
    null;
    r3908 := (r3907);
    r3844 := (r3846 & r3848 & r3850 & r3852 & r3854 & r3856 & r3858 & r3860 & r3862 & r3864 & r3866 & r3868 & r3870 & r3872 & r3874 & r3876 & r3878 & r3880 & r3882 & r3884 & r3886 & r3888 & r3890 & r3892 & r3894 & r3896 & r3898 & r3900 & r3902 & r3904 & r3906 & r3908);
    return r3844;
  end rewire_MetaprogrammingRWw9bdc06a7_3843;
  function rewire_MetaprogrammingRWw80deb1fe_3774 return std_logic_vector
  is
    variable r3839 : std_logic_vector(0 to 0) := (others => '0');
    variable r3838 : std_logic_vector(0 to 0) := (others => '0');
    variable r3837 : std_logic_vector(0 to 0) := (others => '0');
    variable r3836 : std_logic_vector(0 to 0) := (others => '0');
    variable r3835 : std_logic_vector(0 to 0) := (others => '0');
    variable r3834 : std_logic_vector(0 to 0) := (others => '0');
    variable r3833 : std_logic_vector(0 to 0) := (others => '0');
    variable r3832 : std_logic_vector(0 to 0) := (others => '0');
    variable r3831 : std_logic_vector(0 to 0) := (others => '0');
    variable r3830 : std_logic_vector(0 to 0) := (others => '0');
    variable r3829 : std_logic_vector(0 to 0) := (others => '0');
    variable r3828 : std_logic_vector(0 to 0) := (others => '0');
    variable r3827 : std_logic_vector(0 to 0) := (others => '0');
    variable r3826 : std_logic_vector(0 to 0) := (others => '0');
    variable r3825 : std_logic_vector(0 to 0) := (others => '0');
    variable r3824 : std_logic_vector(0 to 0) := (others => '0');
    variable r3823 : std_logic_vector(0 to 0) := (others => '0');
    variable r3822 : std_logic_vector(0 to 0) := (others => '0');
    variable r3821 : std_logic_vector(0 to 0) := (others => '0');
    variable r3820 : std_logic_vector(0 to 0) := (others => '0');
    variable r3819 : std_logic_vector(0 to 0) := (others => '0');
    variable r3818 : std_logic_vector(0 to 0) := (others => '0');
    variable r3817 : std_logic_vector(0 to 0) := (others => '0');
    variable r3816 : std_logic_vector(0 to 0) := (others => '0');
    variable r3815 : std_logic_vector(0 to 0) := (others => '0');
    variable r3814 : std_logic_vector(0 to 0) := (others => '0');
    variable r3813 : std_logic_vector(0 to 0) := (others => '0');
    variable r3812 : std_logic_vector(0 to 0) := (others => '0');
    variable r3811 : std_logic_vector(0 to 0) := (others => '0');
    variable r3810 : std_logic_vector(0 to 0) := (others => '0');
    variable r3809 : std_logic_vector(0 to 0) := (others => '0');
    variable r3808 : std_logic_vector(0 to 0) := (others => '0');
    variable r3807 : std_logic_vector(0 to 0) := (others => '0');
    variable r3806 : std_logic_vector(0 to 0) := (others => '0');
    variable r3805 : std_logic_vector(0 to 0) := (others => '0');
    variable r3804 : std_logic_vector(0 to 0) := (others => '0');
    variable r3803 : std_logic_vector(0 to 0) := (others => '0');
    variable r3802 : std_logic_vector(0 to 0) := (others => '0');
    variable r3801 : std_logic_vector(0 to 0) := (others => '0');
    variable r3800 : std_logic_vector(0 to 0) := (others => '0');
    variable r3799 : std_logic_vector(0 to 0) := (others => '0');
    variable r3798 : std_logic_vector(0 to 0) := (others => '0');
    variable r3797 : std_logic_vector(0 to 0) := (others => '0');
    variable r3796 : std_logic_vector(0 to 0) := (others => '0');
    variable r3795 : std_logic_vector(0 to 0) := (others => '0');
    variable r3794 : std_logic_vector(0 to 0) := (others => '0');
    variable r3793 : std_logic_vector(0 to 0) := (others => '0');
    variable r3792 : std_logic_vector(0 to 0) := (others => '0');
    variable r3791 : std_logic_vector(0 to 0) := (others => '0');
    variable r3790 : std_logic_vector(0 to 0) := (others => '0');
    variable r3789 : std_logic_vector(0 to 0) := (others => '0');
    variable r3788 : std_logic_vector(0 to 0) := (others => '0');
    variable r3787 : std_logic_vector(0 to 0) := (others => '0');
    variable r3786 : std_logic_vector(0 to 0) := (others => '0');
    variable r3785 : std_logic_vector(0 to 0) := (others => '0');
    variable r3784 : std_logic_vector(0 to 0) := (others => '0');
    variable r3783 : std_logic_vector(0 to 0) := (others => '0');
    variable r3782 : std_logic_vector(0 to 0) := (others => '0');
    variable r3781 : std_logic_vector(0 to 0) := (others => '0');
    variable r3780 : std_logic_vector(0 to 0) := (others => '0');
    variable r3779 : std_logic_vector(0 to 0) := (others => '0');
    variable r3778 : std_logic_vector(0 to 0) := (others => '0');
    variable r3777 : std_logic_vector(0 to 0) := (others => '0');
    variable r3776 : std_logic_vector(0 to 0) := (others => '0');
    variable r3775 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r3776 := "1";
    null;
    r3777 := (r3776);
    r3778 := "0";
    null;
    r3779 := (r3778);
    r3780 := "0";
    null;
    r3781 := (r3780);
    r3782 := "0";
    null;
    r3783 := (r3782);
    r3784 := "0";
    null;
    r3785 := (r3784);
    r3786 := "0";
    null;
    r3787 := (r3786);
    r3788 := "0";
    null;
    r3789 := (r3788);
    r3790 := "0";
    null;
    r3791 := (r3790);
    r3792 := "1";
    null;
    r3793 := (r3792);
    r3794 := "1";
    null;
    r3795 := (r3794);
    r3796 := "0";
    null;
    r3797 := (r3796);
    r3798 := "1";
    null;
    r3799 := (r3798);
    r3800 := "1";
    null;
    r3801 := (r3800);
    r3802 := "1";
    null;
    r3803 := (r3802);
    r3804 := "1";
    null;
    r3805 := (r3804);
    r3806 := "0";
    null;
    r3807 := (r3806);
    r3808 := "1";
    null;
    r3809 := (r3808);
    r3810 := "0";
    null;
    r3811 := (r3810);
    r3812 := "1";
    null;
    r3813 := (r3812);
    r3814 := "1";
    null;
    r3815 := (r3814);
    r3816 := "0";
    null;
    r3817 := (r3816);
    r3818 := "0";
    null;
    r3819 := (r3818);
    r3820 := "0";
    null;
    r3821 := (r3820);
    r3822 := "1";
    null;
    r3823 := (r3822);
    r3824 := "1";
    null;
    r3825 := (r3824);
    r3826 := "1";
    null;
    r3827 := (r3826);
    r3828 := "1";
    null;
    r3829 := (r3828);
    r3830 := "1";
    null;
    r3831 := (r3830);
    r3832 := "1";
    null;
    r3833 := (r3832);
    r3834 := "1";
    null;
    r3835 := (r3834);
    r3836 := "1";
    null;
    r3837 := (r3836);
    r3838 := "0";
    null;
    r3839 := (r3838);
    r3775 := (r3777 & r3779 & r3781 & r3783 & r3785 & r3787 & r3789 & r3791 & r3793 & r3795 & r3797 & r3799 & r3801 & r3803 & r3805 & r3807 & r3809 & r3811 & r3813 & r3815 & r3817 & r3819 & r3821 & r3823 & r3825 & r3827 & r3829 & r3831 & r3833 & r3835 & r3837 & r3839);
    return r3775;
  end rewire_MetaprogrammingRWw80deb1fe_3774;
  function rewire_MetaprogrammingRWw72be5d74_3705 return std_logic_vector
  is
    variable r3770 : std_logic_vector(0 to 0) := (others => '0');
    variable r3769 : std_logic_vector(0 to 0) := (others => '0');
    variable r3768 : std_logic_vector(0 to 0) := (others => '0');
    variable r3767 : std_logic_vector(0 to 0) := (others => '0');
    variable r3766 : std_logic_vector(0 to 0) := (others => '0');
    variable r3765 : std_logic_vector(0 to 0) := (others => '0');
    variable r3764 : std_logic_vector(0 to 0) := (others => '0');
    variable r3763 : std_logic_vector(0 to 0) := (others => '0');
    variable r3762 : std_logic_vector(0 to 0) := (others => '0');
    variable r3761 : std_logic_vector(0 to 0) := (others => '0');
    variable r3760 : std_logic_vector(0 to 0) := (others => '0');
    variable r3759 : std_logic_vector(0 to 0) := (others => '0');
    variable r3758 : std_logic_vector(0 to 0) := (others => '0');
    variable r3757 : std_logic_vector(0 to 0) := (others => '0');
    variable r3756 : std_logic_vector(0 to 0) := (others => '0');
    variable r3755 : std_logic_vector(0 to 0) := (others => '0');
    variable r3754 : std_logic_vector(0 to 0) := (others => '0');
    variable r3753 : std_logic_vector(0 to 0) := (others => '0');
    variable r3752 : std_logic_vector(0 to 0) := (others => '0');
    variable r3751 : std_logic_vector(0 to 0) := (others => '0');
    variable r3750 : std_logic_vector(0 to 0) := (others => '0');
    variable r3749 : std_logic_vector(0 to 0) := (others => '0');
    variable r3748 : std_logic_vector(0 to 0) := (others => '0');
    variable r3747 : std_logic_vector(0 to 0) := (others => '0');
    variable r3746 : std_logic_vector(0 to 0) := (others => '0');
    variable r3745 : std_logic_vector(0 to 0) := (others => '0');
    variable r3744 : std_logic_vector(0 to 0) := (others => '0');
    variable r3743 : std_logic_vector(0 to 0) := (others => '0');
    variable r3742 : std_logic_vector(0 to 0) := (others => '0');
    variable r3741 : std_logic_vector(0 to 0) := (others => '0');
    variable r3740 : std_logic_vector(0 to 0) := (others => '0');
    variable r3739 : std_logic_vector(0 to 0) := (others => '0');
    variable r3738 : std_logic_vector(0 to 0) := (others => '0');
    variable r3737 : std_logic_vector(0 to 0) := (others => '0');
    variable r3736 : std_logic_vector(0 to 0) := (others => '0');
    variable r3735 : std_logic_vector(0 to 0) := (others => '0');
    variable r3734 : std_logic_vector(0 to 0) := (others => '0');
    variable r3733 : std_logic_vector(0 to 0) := (others => '0');
    variable r3732 : std_logic_vector(0 to 0) := (others => '0');
    variable r3731 : std_logic_vector(0 to 0) := (others => '0');
    variable r3730 : std_logic_vector(0 to 0) := (others => '0');
    variable r3729 : std_logic_vector(0 to 0) := (others => '0');
    variable r3728 : std_logic_vector(0 to 0) := (others => '0');
    variable r3727 : std_logic_vector(0 to 0) := (others => '0');
    variable r3726 : std_logic_vector(0 to 0) := (others => '0');
    variable r3725 : std_logic_vector(0 to 0) := (others => '0');
    variable r3724 : std_logic_vector(0 to 0) := (others => '0');
    variable r3723 : std_logic_vector(0 to 0) := (others => '0');
    variable r3722 : std_logic_vector(0 to 0) := (others => '0');
    variable r3721 : std_logic_vector(0 to 0) := (others => '0');
    variable r3720 : std_logic_vector(0 to 0) := (others => '0');
    variable r3719 : std_logic_vector(0 to 0) := (others => '0');
    variable r3718 : std_logic_vector(0 to 0) := (others => '0');
    variable r3717 : std_logic_vector(0 to 0) := (others => '0');
    variable r3716 : std_logic_vector(0 to 0) := (others => '0');
    variable r3715 : std_logic_vector(0 to 0) := (others => '0');
    variable r3714 : std_logic_vector(0 to 0) := (others => '0');
    variable r3713 : std_logic_vector(0 to 0) := (others => '0');
    variable r3712 : std_logic_vector(0 to 0) := (others => '0');
    variable r3711 : std_logic_vector(0 to 0) := (others => '0');
    variable r3710 : std_logic_vector(0 to 0) := (others => '0');
    variable r3709 : std_logic_vector(0 to 0) := (others => '0');
    variable r3708 : std_logic_vector(0 to 0) := (others => '0');
    variable r3707 : std_logic_vector(0 to 0) := (others => '0');
    variable r3706 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r3707 := "0";
    null;
    r3708 := (r3707);
    r3709 := "1";
    null;
    r3710 := (r3709);
    r3711 := "1";
    null;
    r3712 := (r3711);
    r3713 := "1";
    null;
    r3714 := (r3713);
    r3715 := "0";
    null;
    r3716 := (r3715);
    r3717 := "0";
    null;
    r3718 := (r3717);
    r3719 := "1";
    null;
    r3720 := (r3719);
    r3721 := "0";
    null;
    r3722 := (r3721);
    r3723 := "1";
    null;
    r3724 := (r3723);
    r3725 := "0";
    null;
    r3726 := (r3725);
    r3727 := "1";
    null;
    r3728 := (r3727);
    r3729 := "1";
    null;
    r3730 := (r3729);
    r3731 := "1";
    null;
    r3732 := (r3731);
    r3733 := "1";
    null;
    r3734 := (r3733);
    r3735 := "1";
    null;
    r3736 := (r3735);
    r3737 := "0";
    null;
    r3738 := (r3737);
    r3739 := "0";
    null;
    r3740 := (r3739);
    r3741 := "1";
    null;
    r3742 := (r3741);
    r3743 := "0";
    null;
    r3744 := (r3743);
    r3745 := "1";
    null;
    r3746 := (r3745);
    r3747 := "1";
    null;
    r3748 := (r3747);
    r3749 := "1";
    null;
    r3750 := (r3749);
    r3751 := "0";
    null;
    r3752 := (r3751);
    r3753 := "1";
    null;
    r3754 := (r3753);
    r3755 := "0";
    null;
    r3756 := (r3755);
    r3757 := "1";
    null;
    r3758 := (r3757);
    r3759 := "1";
    null;
    r3760 := (r3759);
    r3761 := "1";
    null;
    r3762 := (r3761);
    r3763 := "0";
    null;
    r3764 := (r3763);
    r3765 := "1";
    null;
    r3766 := (r3765);
    r3767 := "0";
    null;
    r3768 := (r3767);
    r3769 := "0";
    null;
    r3770 := (r3769);
    r3706 := (r3708 & r3710 & r3712 & r3714 & r3716 & r3718 & r3720 & r3722 & r3724 & r3726 & r3728 & r3730 & r3732 & r3734 & r3736 & r3738 & r3740 & r3742 & r3744 & r3746 & r3748 & r3750 & r3752 & r3754 & r3756 & r3758 & r3760 & r3762 & r3764 & r3766 & r3768 & r3770);
    return r3706;
  end rewire_MetaprogrammingRWw72be5d74_3705;
  function rewire_MetaprogrammingRWw550c7dc3_3636 return std_logic_vector
  is
    variable r3701 : std_logic_vector(0 to 0) := (others => '0');
    variable r3700 : std_logic_vector(0 to 0) := (others => '0');
    variable r3699 : std_logic_vector(0 to 0) := (others => '0');
    variable r3698 : std_logic_vector(0 to 0) := (others => '0');
    variable r3697 : std_logic_vector(0 to 0) := (others => '0');
    variable r3696 : std_logic_vector(0 to 0) := (others => '0');
    variable r3695 : std_logic_vector(0 to 0) := (others => '0');
    variable r3694 : std_logic_vector(0 to 0) := (others => '0');
    variable r3693 : std_logic_vector(0 to 0) := (others => '0');
    variable r3692 : std_logic_vector(0 to 0) := (others => '0');
    variable r3691 : std_logic_vector(0 to 0) := (others => '0');
    variable r3690 : std_logic_vector(0 to 0) := (others => '0');
    variable r3689 : std_logic_vector(0 to 0) := (others => '0');
    variable r3688 : std_logic_vector(0 to 0) := (others => '0');
    variable r3687 : std_logic_vector(0 to 0) := (others => '0');
    variable r3686 : std_logic_vector(0 to 0) := (others => '0');
    variable r3685 : std_logic_vector(0 to 0) := (others => '0');
    variable r3684 : std_logic_vector(0 to 0) := (others => '0');
    variable r3683 : std_logic_vector(0 to 0) := (others => '0');
    variable r3682 : std_logic_vector(0 to 0) := (others => '0');
    variable r3681 : std_logic_vector(0 to 0) := (others => '0');
    variable r3680 : std_logic_vector(0 to 0) := (others => '0');
    variable r3679 : std_logic_vector(0 to 0) := (others => '0');
    variable r3678 : std_logic_vector(0 to 0) := (others => '0');
    variable r3677 : std_logic_vector(0 to 0) := (others => '0');
    variable r3676 : std_logic_vector(0 to 0) := (others => '0');
    variable r3675 : std_logic_vector(0 to 0) := (others => '0');
    variable r3674 : std_logic_vector(0 to 0) := (others => '0');
    variable r3673 : std_logic_vector(0 to 0) := (others => '0');
    variable r3672 : std_logic_vector(0 to 0) := (others => '0');
    variable r3671 : std_logic_vector(0 to 0) := (others => '0');
    variable r3670 : std_logic_vector(0 to 0) := (others => '0');
    variable r3669 : std_logic_vector(0 to 0) := (others => '0');
    variable r3668 : std_logic_vector(0 to 0) := (others => '0');
    variable r3667 : std_logic_vector(0 to 0) := (others => '0');
    variable r3666 : std_logic_vector(0 to 0) := (others => '0');
    variable r3665 : std_logic_vector(0 to 0) := (others => '0');
    variable r3664 : std_logic_vector(0 to 0) := (others => '0');
    variable r3663 : std_logic_vector(0 to 0) := (others => '0');
    variable r3662 : std_logic_vector(0 to 0) := (others => '0');
    variable r3661 : std_logic_vector(0 to 0) := (others => '0');
    variable r3660 : std_logic_vector(0 to 0) := (others => '0');
    variable r3659 : std_logic_vector(0 to 0) := (others => '0');
    variable r3658 : std_logic_vector(0 to 0) := (others => '0');
    variable r3657 : std_logic_vector(0 to 0) := (others => '0');
    variable r3656 : std_logic_vector(0 to 0) := (others => '0');
    variable r3655 : std_logic_vector(0 to 0) := (others => '0');
    variable r3654 : std_logic_vector(0 to 0) := (others => '0');
    variable r3653 : std_logic_vector(0 to 0) := (others => '0');
    variable r3652 : std_logic_vector(0 to 0) := (others => '0');
    variable r3651 : std_logic_vector(0 to 0) := (others => '0');
    variable r3650 : std_logic_vector(0 to 0) := (others => '0');
    variable r3649 : std_logic_vector(0 to 0) := (others => '0');
    variable r3648 : std_logic_vector(0 to 0) := (others => '0');
    variable r3647 : std_logic_vector(0 to 0) := (others => '0');
    variable r3646 : std_logic_vector(0 to 0) := (others => '0');
    variable r3645 : std_logic_vector(0 to 0) := (others => '0');
    variable r3644 : std_logic_vector(0 to 0) := (others => '0');
    variable r3643 : std_logic_vector(0 to 0) := (others => '0');
    variable r3642 : std_logic_vector(0 to 0) := (others => '0');
    variable r3641 : std_logic_vector(0 to 0) := (others => '0');
    variable r3640 : std_logic_vector(0 to 0) := (others => '0');
    variable r3639 : std_logic_vector(0 to 0) := (others => '0');
    variable r3638 : std_logic_vector(0 to 0) := (others => '0');
    variable r3637 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r3638 := "0";
    null;
    r3639 := (r3638);
    r3640 := "1";
    null;
    r3641 := (r3640);
    r3642 := "0";
    null;
    r3643 := (r3642);
    r3644 := "1";
    null;
    r3645 := (r3644);
    r3646 := "0";
    null;
    r3647 := (r3646);
    r3648 := "1";
    null;
    r3649 := (r3648);
    r3650 := "0";
    null;
    r3651 := (r3650);
    r3652 := "1";
    null;
    r3653 := (r3652);
    r3654 := "0";
    null;
    r3655 := (r3654);
    r3656 := "0";
    null;
    r3657 := (r3656);
    r3658 := "0";
    null;
    r3659 := (r3658);
    r3660 := "0";
    null;
    r3661 := (r3660);
    r3662 := "1";
    null;
    r3663 := (r3662);
    r3664 := "1";
    null;
    r3665 := (r3664);
    r3666 := "0";
    null;
    r3667 := (r3666);
    r3668 := "0";
    null;
    r3669 := (r3668);
    r3670 := "0";
    null;
    r3671 := (r3670);
    r3672 := "1";
    null;
    r3673 := (r3672);
    r3674 := "1";
    null;
    r3675 := (r3674);
    r3676 := "1";
    null;
    r3677 := (r3676);
    r3678 := "1";
    null;
    r3679 := (r3678);
    r3680 := "1";
    null;
    r3681 := (r3680);
    r3682 := "0";
    null;
    r3683 := (r3682);
    r3684 := "1";
    null;
    r3685 := (r3684);
    r3686 := "1";
    null;
    r3687 := (r3686);
    r3688 := "1";
    null;
    r3689 := (r3688);
    r3690 := "0";
    null;
    r3691 := (r3690);
    r3692 := "0";
    null;
    r3693 := (r3692);
    r3694 := "0";
    null;
    r3695 := (r3694);
    r3696 := "0";
    null;
    r3697 := (r3696);
    r3698 := "1";
    null;
    r3699 := (r3698);
    r3700 := "1";
    null;
    r3701 := (r3700);
    r3637 := (r3639 & r3641 & r3643 & r3645 & r3647 & r3649 & r3651 & r3653 & r3655 & r3657 & r3659 & r3661 & r3663 & r3665 & r3667 & r3669 & r3671 & r3673 & r3675 & r3677 & r3679 & r3681 & r3683 & r3685 & r3687 & r3689 & r3691 & r3693 & r3695 & r3697 & r3699 & r3701);
    return r3637;
  end rewire_MetaprogrammingRWw550c7dc3_3636;
  function rewire_MetaprogrammingRWw243185be_3567 return std_logic_vector
  is
    variable r3632 : std_logic_vector(0 to 0) := (others => '0');
    variable r3631 : std_logic_vector(0 to 0) := (others => '0');
    variable r3630 : std_logic_vector(0 to 0) := (others => '0');
    variable r3629 : std_logic_vector(0 to 0) := (others => '0');
    variable r3628 : std_logic_vector(0 to 0) := (others => '0');
    variable r3627 : std_logic_vector(0 to 0) := (others => '0');
    variable r3626 : std_logic_vector(0 to 0) := (others => '0');
    variable r3625 : std_logic_vector(0 to 0) := (others => '0');
    variable r3624 : std_logic_vector(0 to 0) := (others => '0');
    variable r3623 : std_logic_vector(0 to 0) := (others => '0');
    variable r3622 : std_logic_vector(0 to 0) := (others => '0');
    variable r3621 : std_logic_vector(0 to 0) := (others => '0');
    variable r3620 : std_logic_vector(0 to 0) := (others => '0');
    variable r3619 : std_logic_vector(0 to 0) := (others => '0');
    variable r3618 : std_logic_vector(0 to 0) := (others => '0');
    variable r3617 : std_logic_vector(0 to 0) := (others => '0');
    variable r3616 : std_logic_vector(0 to 0) := (others => '0');
    variable r3615 : std_logic_vector(0 to 0) := (others => '0');
    variable r3614 : std_logic_vector(0 to 0) := (others => '0');
    variable r3613 : std_logic_vector(0 to 0) := (others => '0');
    variable r3612 : std_logic_vector(0 to 0) := (others => '0');
    variable r3611 : std_logic_vector(0 to 0) := (others => '0');
    variable r3610 : std_logic_vector(0 to 0) := (others => '0');
    variable r3609 : std_logic_vector(0 to 0) := (others => '0');
    variable r3608 : std_logic_vector(0 to 0) := (others => '0');
    variable r3607 : std_logic_vector(0 to 0) := (others => '0');
    variable r3606 : std_logic_vector(0 to 0) := (others => '0');
    variable r3605 : std_logic_vector(0 to 0) := (others => '0');
    variable r3604 : std_logic_vector(0 to 0) := (others => '0');
    variable r3603 : std_logic_vector(0 to 0) := (others => '0');
    variable r3602 : std_logic_vector(0 to 0) := (others => '0');
    variable r3601 : std_logic_vector(0 to 0) := (others => '0');
    variable r3600 : std_logic_vector(0 to 0) := (others => '0');
    variable r3599 : std_logic_vector(0 to 0) := (others => '0');
    variable r3598 : std_logic_vector(0 to 0) := (others => '0');
    variable r3597 : std_logic_vector(0 to 0) := (others => '0');
    variable r3596 : std_logic_vector(0 to 0) := (others => '0');
    variable r3595 : std_logic_vector(0 to 0) := (others => '0');
    variable r3594 : std_logic_vector(0 to 0) := (others => '0');
    variable r3593 : std_logic_vector(0 to 0) := (others => '0');
    variable r3592 : std_logic_vector(0 to 0) := (others => '0');
    variable r3591 : std_logic_vector(0 to 0) := (others => '0');
    variable r3590 : std_logic_vector(0 to 0) := (others => '0');
    variable r3589 : std_logic_vector(0 to 0) := (others => '0');
    variable r3588 : std_logic_vector(0 to 0) := (others => '0');
    variable r3587 : std_logic_vector(0 to 0) := (others => '0');
    variable r3586 : std_logic_vector(0 to 0) := (others => '0');
    variable r3585 : std_logic_vector(0 to 0) := (others => '0');
    variable r3584 : std_logic_vector(0 to 0) := (others => '0');
    variable r3583 : std_logic_vector(0 to 0) := (others => '0');
    variable r3582 : std_logic_vector(0 to 0) := (others => '0');
    variable r3581 : std_logic_vector(0 to 0) := (others => '0');
    variable r3580 : std_logic_vector(0 to 0) := (others => '0');
    variable r3579 : std_logic_vector(0 to 0) := (others => '0');
    variable r3578 : std_logic_vector(0 to 0) := (others => '0');
    variable r3577 : std_logic_vector(0 to 0) := (others => '0');
    variable r3576 : std_logic_vector(0 to 0) := (others => '0');
    variable r3575 : std_logic_vector(0 to 0) := (others => '0');
    variable r3574 : std_logic_vector(0 to 0) := (others => '0');
    variable r3573 : std_logic_vector(0 to 0) := (others => '0');
    variable r3572 : std_logic_vector(0 to 0) := (others => '0');
    variable r3571 : std_logic_vector(0 to 0) := (others => '0');
    variable r3570 : std_logic_vector(0 to 0) := (others => '0');
    variable r3569 : std_logic_vector(0 to 0) := (others => '0');
    variable r3568 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r3569 := "0";
    null;
    r3570 := (r3569);
    r3571 := "0";
    null;
    r3572 := (r3571);
    r3573 := "1";
    null;
    r3574 := (r3573);
    r3575 := "0";
    null;
    r3576 := (r3575);
    r3577 := "0";
    null;
    r3578 := (r3577);
    r3579 := "1";
    null;
    r3580 := (r3579);
    r3581 := "0";
    null;
    r3582 := (r3581);
    r3583 := "0";
    null;
    r3584 := (r3583);
    r3585 := "0";
    null;
    r3586 := (r3585);
    r3587 := "0";
    null;
    r3588 := (r3587);
    r3589 := "1";
    null;
    r3590 := (r3589);
    r3591 := "1";
    null;
    r3592 := (r3591);
    r3593 := "0";
    null;
    r3594 := (r3593);
    r3595 := "0";
    null;
    r3596 := (r3595);
    r3597 := "0";
    null;
    r3598 := (r3597);
    r3599 := "1";
    null;
    r3600 := (r3599);
    r3601 := "1";
    null;
    r3602 := (r3601);
    r3603 := "0";
    null;
    r3604 := (r3603);
    r3605 := "0";
    null;
    r3606 := (r3605);
    r3607 := "0";
    null;
    r3608 := (r3607);
    r3609 := "0";
    null;
    r3610 := (r3609);
    r3611 := "1";
    null;
    r3612 := (r3611);
    r3613 := "0";
    null;
    r3614 := (r3613);
    r3615 := "1";
    null;
    r3616 := (r3615);
    r3617 := "1";
    null;
    r3618 := (r3617);
    r3619 := "0";
    null;
    r3620 := (r3619);
    r3621 := "1";
    null;
    r3622 := (r3621);
    r3623 := "1";
    null;
    r3624 := (r3623);
    r3625 := "1";
    null;
    r3626 := (r3625);
    r3627 := "1";
    null;
    r3628 := (r3627);
    r3629 := "1";
    null;
    r3630 := (r3629);
    r3631 := "0";
    null;
    r3632 := (r3631);
    r3568 := (r3570 & r3572 & r3574 & r3576 & r3578 & r3580 & r3582 & r3584 & r3586 & r3588 & r3590 & r3592 & r3594 & r3596 & r3598 & r3600 & r3602 & r3604 & r3606 & r3608 & r3610 & r3612 & r3614 & r3616 & r3618 & r3620 & r3622 & r3624 & r3626 & r3628 & r3630 & r3632);
    return r3568;
  end rewire_MetaprogrammingRWw243185be_3567;
  function rewire_MetaprogrammingRWw12835b01_3498 return std_logic_vector
  is
    variable r3563 : std_logic_vector(0 to 0) := (others => '0');
    variable r3562 : std_logic_vector(0 to 0) := (others => '0');
    variable r3561 : std_logic_vector(0 to 0) := (others => '0');
    variable r3560 : std_logic_vector(0 to 0) := (others => '0');
    variable r3559 : std_logic_vector(0 to 0) := (others => '0');
    variable r3558 : std_logic_vector(0 to 0) := (others => '0');
    variable r3557 : std_logic_vector(0 to 0) := (others => '0');
    variable r3556 : std_logic_vector(0 to 0) := (others => '0');
    variable r3555 : std_logic_vector(0 to 0) := (others => '0');
    variable r3554 : std_logic_vector(0 to 0) := (others => '0');
    variable r3553 : std_logic_vector(0 to 0) := (others => '0');
    variable r3552 : std_logic_vector(0 to 0) := (others => '0');
    variable r3551 : std_logic_vector(0 to 0) := (others => '0');
    variable r3550 : std_logic_vector(0 to 0) := (others => '0');
    variable r3549 : std_logic_vector(0 to 0) := (others => '0');
    variable r3548 : std_logic_vector(0 to 0) := (others => '0');
    variable r3547 : std_logic_vector(0 to 0) := (others => '0');
    variable r3546 : std_logic_vector(0 to 0) := (others => '0');
    variable r3545 : std_logic_vector(0 to 0) := (others => '0');
    variable r3544 : std_logic_vector(0 to 0) := (others => '0');
    variable r3543 : std_logic_vector(0 to 0) := (others => '0');
    variable r3542 : std_logic_vector(0 to 0) := (others => '0');
    variable r3541 : std_logic_vector(0 to 0) := (others => '0');
    variable r3540 : std_logic_vector(0 to 0) := (others => '0');
    variable r3539 : std_logic_vector(0 to 0) := (others => '0');
    variable r3538 : std_logic_vector(0 to 0) := (others => '0');
    variable r3537 : std_logic_vector(0 to 0) := (others => '0');
    variable r3536 : std_logic_vector(0 to 0) := (others => '0');
    variable r3535 : std_logic_vector(0 to 0) := (others => '0');
    variable r3534 : std_logic_vector(0 to 0) := (others => '0');
    variable r3533 : std_logic_vector(0 to 0) := (others => '0');
    variable r3532 : std_logic_vector(0 to 0) := (others => '0');
    variable r3531 : std_logic_vector(0 to 0) := (others => '0');
    variable r3530 : std_logic_vector(0 to 0) := (others => '0');
    variable r3529 : std_logic_vector(0 to 0) := (others => '0');
    variable r3528 : std_logic_vector(0 to 0) := (others => '0');
    variable r3527 : std_logic_vector(0 to 0) := (others => '0');
    variable r3526 : std_logic_vector(0 to 0) := (others => '0');
    variable r3525 : std_logic_vector(0 to 0) := (others => '0');
    variable r3524 : std_logic_vector(0 to 0) := (others => '0');
    variable r3523 : std_logic_vector(0 to 0) := (others => '0');
    variable r3522 : std_logic_vector(0 to 0) := (others => '0');
    variable r3521 : std_logic_vector(0 to 0) := (others => '0');
    variable r3520 : std_logic_vector(0 to 0) := (others => '0');
    variable r3519 : std_logic_vector(0 to 0) := (others => '0');
    variable r3518 : std_logic_vector(0 to 0) := (others => '0');
    variable r3517 : std_logic_vector(0 to 0) := (others => '0');
    variable r3516 : std_logic_vector(0 to 0) := (others => '0');
    variable r3515 : std_logic_vector(0 to 0) := (others => '0');
    variable r3514 : std_logic_vector(0 to 0) := (others => '0');
    variable r3513 : std_logic_vector(0 to 0) := (others => '0');
    variable r3512 : std_logic_vector(0 to 0) := (others => '0');
    variable r3511 : std_logic_vector(0 to 0) := (others => '0');
    variable r3510 : std_logic_vector(0 to 0) := (others => '0');
    variable r3509 : std_logic_vector(0 to 0) := (others => '0');
    variable r3508 : std_logic_vector(0 to 0) := (others => '0');
    variable r3507 : std_logic_vector(0 to 0) := (others => '0');
    variable r3506 : std_logic_vector(0 to 0) := (others => '0');
    variable r3505 : std_logic_vector(0 to 0) := (others => '0');
    variable r3504 : std_logic_vector(0 to 0) := (others => '0');
    variable r3503 : std_logic_vector(0 to 0) := (others => '0');
    variable r3502 : std_logic_vector(0 to 0) := (others => '0');
    variable r3501 : std_logic_vector(0 to 0) := (others => '0');
    variable r3500 : std_logic_vector(0 to 0) := (others => '0');
    variable r3499 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r3500 := "0";
    null;
    r3501 := (r3500);
    r3502 := "0";
    null;
    r3503 := (r3502);
    r3504 := "0";
    null;
    r3505 := (r3504);
    r3506 := "1";
    null;
    r3507 := (r3506);
    r3508 := "0";
    null;
    r3509 := (r3508);
    r3510 := "0";
    null;
    r3511 := (r3510);
    r3512 := "1";
    null;
    r3513 := (r3512);
    r3514 := "0";
    null;
    r3515 := (r3514);
    r3516 := "1";
    null;
    r3517 := (r3516);
    r3518 := "0";
    null;
    r3519 := (r3518);
    r3520 := "0";
    null;
    r3521 := (r3520);
    r3522 := "0";
    null;
    r3523 := (r3522);
    r3524 := "0";
    null;
    r3525 := (r3524);
    r3526 := "0";
    null;
    r3527 := (r3526);
    r3528 := "1";
    null;
    r3529 := (r3528);
    r3530 := "1";
    null;
    r3531 := (r3530);
    r3532 := "0";
    null;
    r3533 := (r3532);
    r3534 := "1";
    null;
    r3535 := (r3534);
    r3536 := "0";
    null;
    r3537 := (r3536);
    r3538 := "1";
    null;
    r3539 := (r3538);
    r3540 := "1";
    null;
    r3541 := (r3540);
    r3542 := "0";
    null;
    r3543 := (r3542);
    r3544 := "1";
    null;
    r3545 := (r3544);
    r3546 := "1";
    null;
    r3547 := (r3546);
    r3548 := "0";
    null;
    r3549 := (r3548);
    r3550 := "0";
    null;
    r3551 := (r3550);
    r3552 := "0";
    null;
    r3553 := (r3552);
    r3554 := "0";
    null;
    r3555 := (r3554);
    r3556 := "0";
    null;
    r3557 := (r3556);
    r3558 := "0";
    null;
    r3559 := (r3558);
    r3560 := "0";
    null;
    r3561 := (r3560);
    r3562 := "1";
    null;
    r3563 := (r3562);
    r3499 := (r3501 & r3503 & r3505 & r3507 & r3509 & r3511 & r3513 & r3515 & r3517 & r3519 & r3521 & r3523 & r3525 & r3527 & r3529 & r3531 & r3533 & r3535 & r3537 & r3539 & r3541 & r3543 & r3545 & r3547 & r3549 & r3551 & r3553 & r3555 & r3557 & r3559 & r3561 & r3563);
    return r3499;
  end rewire_MetaprogrammingRWw12835b01_3498;
  function rewire_MetaprogrammingRWwd807aa98_3429 return std_logic_vector
  is
    variable r3494 : std_logic_vector(0 to 0) := (others => '0');
    variable r3493 : std_logic_vector(0 to 0) := (others => '0');
    variable r3492 : std_logic_vector(0 to 0) := (others => '0');
    variable r3491 : std_logic_vector(0 to 0) := (others => '0');
    variable r3490 : std_logic_vector(0 to 0) := (others => '0');
    variable r3489 : std_logic_vector(0 to 0) := (others => '0');
    variable r3488 : std_logic_vector(0 to 0) := (others => '0');
    variable r3487 : std_logic_vector(0 to 0) := (others => '0');
    variable r3486 : std_logic_vector(0 to 0) := (others => '0');
    variable r3485 : std_logic_vector(0 to 0) := (others => '0');
    variable r3484 : std_logic_vector(0 to 0) := (others => '0');
    variable r3483 : std_logic_vector(0 to 0) := (others => '0');
    variable r3482 : std_logic_vector(0 to 0) := (others => '0');
    variable r3481 : std_logic_vector(0 to 0) := (others => '0');
    variable r3480 : std_logic_vector(0 to 0) := (others => '0');
    variable r3479 : std_logic_vector(0 to 0) := (others => '0');
    variable r3478 : std_logic_vector(0 to 0) := (others => '0');
    variable r3477 : std_logic_vector(0 to 0) := (others => '0');
    variable r3476 : std_logic_vector(0 to 0) := (others => '0');
    variable r3475 : std_logic_vector(0 to 0) := (others => '0');
    variable r3474 : std_logic_vector(0 to 0) := (others => '0');
    variable r3473 : std_logic_vector(0 to 0) := (others => '0');
    variable r3472 : std_logic_vector(0 to 0) := (others => '0');
    variable r3471 : std_logic_vector(0 to 0) := (others => '0');
    variable r3470 : std_logic_vector(0 to 0) := (others => '0');
    variable r3469 : std_logic_vector(0 to 0) := (others => '0');
    variable r3468 : std_logic_vector(0 to 0) := (others => '0');
    variable r3467 : std_logic_vector(0 to 0) := (others => '0');
    variable r3466 : std_logic_vector(0 to 0) := (others => '0');
    variable r3465 : std_logic_vector(0 to 0) := (others => '0');
    variable r3464 : std_logic_vector(0 to 0) := (others => '0');
    variable r3463 : std_logic_vector(0 to 0) := (others => '0');
    variable r3462 : std_logic_vector(0 to 0) := (others => '0');
    variable r3461 : std_logic_vector(0 to 0) := (others => '0');
    variable r3460 : std_logic_vector(0 to 0) := (others => '0');
    variable r3459 : std_logic_vector(0 to 0) := (others => '0');
    variable r3458 : std_logic_vector(0 to 0) := (others => '0');
    variable r3457 : std_logic_vector(0 to 0) := (others => '0');
    variable r3456 : std_logic_vector(0 to 0) := (others => '0');
    variable r3455 : std_logic_vector(0 to 0) := (others => '0');
    variable r3454 : std_logic_vector(0 to 0) := (others => '0');
    variable r3453 : std_logic_vector(0 to 0) := (others => '0');
    variable r3452 : std_logic_vector(0 to 0) := (others => '0');
    variable r3451 : std_logic_vector(0 to 0) := (others => '0');
    variable r3450 : std_logic_vector(0 to 0) := (others => '0');
    variable r3449 : std_logic_vector(0 to 0) := (others => '0');
    variable r3448 : std_logic_vector(0 to 0) := (others => '0');
    variable r3447 : std_logic_vector(0 to 0) := (others => '0');
    variable r3446 : std_logic_vector(0 to 0) := (others => '0');
    variable r3445 : std_logic_vector(0 to 0) := (others => '0');
    variable r3444 : std_logic_vector(0 to 0) := (others => '0');
    variable r3443 : std_logic_vector(0 to 0) := (others => '0');
    variable r3442 : std_logic_vector(0 to 0) := (others => '0');
    variable r3441 : std_logic_vector(0 to 0) := (others => '0');
    variable r3440 : std_logic_vector(0 to 0) := (others => '0');
    variable r3439 : std_logic_vector(0 to 0) := (others => '0');
    variable r3438 : std_logic_vector(0 to 0) := (others => '0');
    variable r3437 : std_logic_vector(0 to 0) := (others => '0');
    variable r3436 : std_logic_vector(0 to 0) := (others => '0');
    variable r3435 : std_logic_vector(0 to 0) := (others => '0');
    variable r3434 : std_logic_vector(0 to 0) := (others => '0');
    variable r3433 : std_logic_vector(0 to 0) := (others => '0');
    variable r3432 : std_logic_vector(0 to 0) := (others => '0');
    variable r3431 : std_logic_vector(0 to 0) := (others => '0');
    variable r3430 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r3431 := "1";
    null;
    r3432 := (r3431);
    r3433 := "1";
    null;
    r3434 := (r3433);
    r3435 := "0";
    null;
    r3436 := (r3435);
    r3437 := "1";
    null;
    r3438 := (r3437);
    r3439 := "1";
    null;
    r3440 := (r3439);
    r3441 := "0";
    null;
    r3442 := (r3441);
    r3443 := "0";
    null;
    r3444 := (r3443);
    r3445 := "0";
    null;
    r3446 := (r3445);
    r3447 := "0";
    null;
    r3448 := (r3447);
    r3449 := "0";
    null;
    r3450 := (r3449);
    r3451 := "0";
    null;
    r3452 := (r3451);
    r3453 := "0";
    null;
    r3454 := (r3453);
    r3455 := "0";
    null;
    r3456 := (r3455);
    r3457 := "1";
    null;
    r3458 := (r3457);
    r3459 := "1";
    null;
    r3460 := (r3459);
    r3461 := "1";
    null;
    r3462 := (r3461);
    r3463 := "1";
    null;
    r3464 := (r3463);
    r3465 := "0";
    null;
    r3466 := (r3465);
    r3467 := "1";
    null;
    r3468 := (r3467);
    r3469 := "0";
    null;
    r3470 := (r3469);
    r3471 := "1";
    null;
    r3472 := (r3471);
    r3473 := "0";
    null;
    r3474 := (r3473);
    r3475 := "1";
    null;
    r3476 := (r3475);
    r3477 := "0";
    null;
    r3478 := (r3477);
    r3479 := "1";
    null;
    r3480 := (r3479);
    r3481 := "0";
    null;
    r3482 := (r3481);
    r3483 := "0";
    null;
    r3484 := (r3483);
    r3485 := "1";
    null;
    r3486 := (r3485);
    r3487 := "1";
    null;
    r3488 := (r3487);
    r3489 := "0";
    null;
    r3490 := (r3489);
    r3491 := "0";
    null;
    r3492 := (r3491);
    r3493 := "0";
    null;
    r3494 := (r3493);
    r3430 := (r3432 & r3434 & r3436 & r3438 & r3440 & r3442 & r3444 & r3446 & r3448 & r3450 & r3452 & r3454 & r3456 & r3458 & r3460 & r3462 & r3464 & r3466 & r3468 & r3470 & r3472 & r3474 & r3476 & r3478 & r3480 & r3482 & r3484 & r3486 & r3488 & r3490 & r3492 & r3494);
    return r3430;
  end rewire_MetaprogrammingRWwd807aa98_3429;
  function rewire_MetaprogrammingRWwab1c5ed5_3360 return std_logic_vector
  is
    variable r3425 : std_logic_vector(0 to 0) := (others => '0');
    variable r3424 : std_logic_vector(0 to 0) := (others => '0');
    variable r3423 : std_logic_vector(0 to 0) := (others => '0');
    variable r3422 : std_logic_vector(0 to 0) := (others => '0');
    variable r3421 : std_logic_vector(0 to 0) := (others => '0');
    variable r3420 : std_logic_vector(0 to 0) := (others => '0');
    variable r3419 : std_logic_vector(0 to 0) := (others => '0');
    variable r3418 : std_logic_vector(0 to 0) := (others => '0');
    variable r3417 : std_logic_vector(0 to 0) := (others => '0');
    variable r3416 : std_logic_vector(0 to 0) := (others => '0');
    variable r3415 : std_logic_vector(0 to 0) := (others => '0');
    variable r3414 : std_logic_vector(0 to 0) := (others => '0');
    variable r3413 : std_logic_vector(0 to 0) := (others => '0');
    variable r3412 : std_logic_vector(0 to 0) := (others => '0');
    variable r3411 : std_logic_vector(0 to 0) := (others => '0');
    variable r3410 : std_logic_vector(0 to 0) := (others => '0');
    variable r3409 : std_logic_vector(0 to 0) := (others => '0');
    variable r3408 : std_logic_vector(0 to 0) := (others => '0');
    variable r3407 : std_logic_vector(0 to 0) := (others => '0');
    variable r3406 : std_logic_vector(0 to 0) := (others => '0');
    variable r3405 : std_logic_vector(0 to 0) := (others => '0');
    variable r3404 : std_logic_vector(0 to 0) := (others => '0');
    variable r3403 : std_logic_vector(0 to 0) := (others => '0');
    variable r3402 : std_logic_vector(0 to 0) := (others => '0');
    variable r3401 : std_logic_vector(0 to 0) := (others => '0');
    variable r3400 : std_logic_vector(0 to 0) := (others => '0');
    variable r3399 : std_logic_vector(0 to 0) := (others => '0');
    variable r3398 : std_logic_vector(0 to 0) := (others => '0');
    variable r3397 : std_logic_vector(0 to 0) := (others => '0');
    variable r3396 : std_logic_vector(0 to 0) := (others => '0');
    variable r3395 : std_logic_vector(0 to 0) := (others => '0');
    variable r3394 : std_logic_vector(0 to 0) := (others => '0');
    variable r3393 : std_logic_vector(0 to 0) := (others => '0');
    variable r3392 : std_logic_vector(0 to 0) := (others => '0');
    variable r3391 : std_logic_vector(0 to 0) := (others => '0');
    variable r3390 : std_logic_vector(0 to 0) := (others => '0');
    variable r3389 : std_logic_vector(0 to 0) := (others => '0');
    variable r3388 : std_logic_vector(0 to 0) := (others => '0');
    variable r3387 : std_logic_vector(0 to 0) := (others => '0');
    variable r3386 : std_logic_vector(0 to 0) := (others => '0');
    variable r3385 : std_logic_vector(0 to 0) := (others => '0');
    variable r3384 : std_logic_vector(0 to 0) := (others => '0');
    variable r3383 : std_logic_vector(0 to 0) := (others => '0');
    variable r3382 : std_logic_vector(0 to 0) := (others => '0');
    variable r3381 : std_logic_vector(0 to 0) := (others => '0');
    variable r3380 : std_logic_vector(0 to 0) := (others => '0');
    variable r3379 : std_logic_vector(0 to 0) := (others => '0');
    variable r3378 : std_logic_vector(0 to 0) := (others => '0');
    variable r3377 : std_logic_vector(0 to 0) := (others => '0');
    variable r3376 : std_logic_vector(0 to 0) := (others => '0');
    variable r3375 : std_logic_vector(0 to 0) := (others => '0');
    variable r3374 : std_logic_vector(0 to 0) := (others => '0');
    variable r3373 : std_logic_vector(0 to 0) := (others => '0');
    variable r3372 : std_logic_vector(0 to 0) := (others => '0');
    variable r3371 : std_logic_vector(0 to 0) := (others => '0');
    variable r3370 : std_logic_vector(0 to 0) := (others => '0');
    variable r3369 : std_logic_vector(0 to 0) := (others => '0');
    variable r3368 : std_logic_vector(0 to 0) := (others => '0');
    variable r3367 : std_logic_vector(0 to 0) := (others => '0');
    variable r3366 : std_logic_vector(0 to 0) := (others => '0');
    variable r3365 : std_logic_vector(0 to 0) := (others => '0');
    variable r3364 : std_logic_vector(0 to 0) := (others => '0');
    variable r3363 : std_logic_vector(0 to 0) := (others => '0');
    variable r3362 : std_logic_vector(0 to 0) := (others => '0');
    variable r3361 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r3362 := "1";
    null;
    r3363 := (r3362);
    r3364 := "0";
    null;
    r3365 := (r3364);
    r3366 := "1";
    null;
    r3367 := (r3366);
    r3368 := "0";
    null;
    r3369 := (r3368);
    r3370 := "1";
    null;
    r3371 := (r3370);
    r3372 := "0";
    null;
    r3373 := (r3372);
    r3374 := "1";
    null;
    r3375 := (r3374);
    r3376 := "1";
    null;
    r3377 := (r3376);
    r3378 := "0";
    null;
    r3379 := (r3378);
    r3380 := "0";
    null;
    r3381 := (r3380);
    r3382 := "0";
    null;
    r3383 := (r3382);
    r3384 := "1";
    null;
    r3385 := (r3384);
    r3386 := "1";
    null;
    r3387 := (r3386);
    r3388 := "1";
    null;
    r3389 := (r3388);
    r3390 := "0";
    null;
    r3391 := (r3390);
    r3392 := "0";
    null;
    r3393 := (r3392);
    r3394 := "0";
    null;
    r3395 := (r3394);
    r3396 := "1";
    null;
    r3397 := (r3396);
    r3398 := "0";
    null;
    r3399 := (r3398);
    r3400 := "1";
    null;
    r3401 := (r3400);
    r3402 := "1";
    null;
    r3403 := (r3402);
    r3404 := "1";
    null;
    r3405 := (r3404);
    r3406 := "1";
    null;
    r3407 := (r3406);
    r3408 := "0";
    null;
    r3409 := (r3408);
    r3410 := "1";
    null;
    r3411 := (r3410);
    r3412 := "1";
    null;
    r3413 := (r3412);
    r3414 := "0";
    null;
    r3415 := (r3414);
    r3416 := "1";
    null;
    r3417 := (r3416);
    r3418 := "0";
    null;
    r3419 := (r3418);
    r3420 := "1";
    null;
    r3421 := (r3420);
    r3422 := "0";
    null;
    r3423 := (r3422);
    r3424 := "1";
    null;
    r3425 := (r3424);
    r3361 := (r3363 & r3365 & r3367 & r3369 & r3371 & r3373 & r3375 & r3377 & r3379 & r3381 & r3383 & r3385 & r3387 & r3389 & r3391 & r3393 & r3395 & r3397 & r3399 & r3401 & r3403 & r3405 & r3407 & r3409 & r3411 & r3413 & r3415 & r3417 & r3419 & r3421 & r3423 & r3425);
    return r3361;
  end rewire_MetaprogrammingRWwab1c5ed5_3360;
  function rewire_MetaprogrammingRWw923f82a4_3291 return std_logic_vector
  is
    variable r3356 : std_logic_vector(0 to 0) := (others => '0');
    variable r3355 : std_logic_vector(0 to 0) := (others => '0');
    variable r3354 : std_logic_vector(0 to 0) := (others => '0');
    variable r3353 : std_logic_vector(0 to 0) := (others => '0');
    variable r3352 : std_logic_vector(0 to 0) := (others => '0');
    variable r3351 : std_logic_vector(0 to 0) := (others => '0');
    variable r3350 : std_logic_vector(0 to 0) := (others => '0');
    variable r3349 : std_logic_vector(0 to 0) := (others => '0');
    variable r3348 : std_logic_vector(0 to 0) := (others => '0');
    variable r3347 : std_logic_vector(0 to 0) := (others => '0');
    variable r3346 : std_logic_vector(0 to 0) := (others => '0');
    variable r3345 : std_logic_vector(0 to 0) := (others => '0');
    variable r3344 : std_logic_vector(0 to 0) := (others => '0');
    variable r3343 : std_logic_vector(0 to 0) := (others => '0');
    variable r3342 : std_logic_vector(0 to 0) := (others => '0');
    variable r3341 : std_logic_vector(0 to 0) := (others => '0');
    variable r3340 : std_logic_vector(0 to 0) := (others => '0');
    variable r3339 : std_logic_vector(0 to 0) := (others => '0');
    variable r3338 : std_logic_vector(0 to 0) := (others => '0');
    variable r3337 : std_logic_vector(0 to 0) := (others => '0');
    variable r3336 : std_logic_vector(0 to 0) := (others => '0');
    variable r3335 : std_logic_vector(0 to 0) := (others => '0');
    variable r3334 : std_logic_vector(0 to 0) := (others => '0');
    variable r3333 : std_logic_vector(0 to 0) := (others => '0');
    variable r3332 : std_logic_vector(0 to 0) := (others => '0');
    variable r3331 : std_logic_vector(0 to 0) := (others => '0');
    variable r3330 : std_logic_vector(0 to 0) := (others => '0');
    variable r3329 : std_logic_vector(0 to 0) := (others => '0');
    variable r3328 : std_logic_vector(0 to 0) := (others => '0');
    variable r3327 : std_logic_vector(0 to 0) := (others => '0');
    variable r3326 : std_logic_vector(0 to 0) := (others => '0');
    variable r3325 : std_logic_vector(0 to 0) := (others => '0');
    variable r3324 : std_logic_vector(0 to 0) := (others => '0');
    variable r3323 : std_logic_vector(0 to 0) := (others => '0');
    variable r3322 : std_logic_vector(0 to 0) := (others => '0');
    variable r3321 : std_logic_vector(0 to 0) := (others => '0');
    variable r3320 : std_logic_vector(0 to 0) := (others => '0');
    variable r3319 : std_logic_vector(0 to 0) := (others => '0');
    variable r3318 : std_logic_vector(0 to 0) := (others => '0');
    variable r3317 : std_logic_vector(0 to 0) := (others => '0');
    variable r3316 : std_logic_vector(0 to 0) := (others => '0');
    variable r3315 : std_logic_vector(0 to 0) := (others => '0');
    variable r3314 : std_logic_vector(0 to 0) := (others => '0');
    variable r3313 : std_logic_vector(0 to 0) := (others => '0');
    variable r3312 : std_logic_vector(0 to 0) := (others => '0');
    variable r3311 : std_logic_vector(0 to 0) := (others => '0');
    variable r3310 : std_logic_vector(0 to 0) := (others => '0');
    variable r3309 : std_logic_vector(0 to 0) := (others => '0');
    variable r3308 : std_logic_vector(0 to 0) := (others => '0');
    variable r3307 : std_logic_vector(0 to 0) := (others => '0');
    variable r3306 : std_logic_vector(0 to 0) := (others => '0');
    variable r3305 : std_logic_vector(0 to 0) := (others => '0');
    variable r3304 : std_logic_vector(0 to 0) := (others => '0');
    variable r3303 : std_logic_vector(0 to 0) := (others => '0');
    variable r3302 : std_logic_vector(0 to 0) := (others => '0');
    variable r3301 : std_logic_vector(0 to 0) := (others => '0');
    variable r3300 : std_logic_vector(0 to 0) := (others => '0');
    variable r3299 : std_logic_vector(0 to 0) := (others => '0');
    variable r3298 : std_logic_vector(0 to 0) := (others => '0');
    variable r3297 : std_logic_vector(0 to 0) := (others => '0');
    variable r3296 : std_logic_vector(0 to 0) := (others => '0');
    variable r3295 : std_logic_vector(0 to 0) := (others => '0');
    variable r3294 : std_logic_vector(0 to 0) := (others => '0');
    variable r3293 : std_logic_vector(0 to 0) := (others => '0');
    variable r3292 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r3293 := "1";
    null;
    r3294 := (r3293);
    r3295 := "0";
    null;
    r3296 := (r3295);
    r3297 := "0";
    null;
    r3298 := (r3297);
    r3299 := "1";
    null;
    r3300 := (r3299);
    r3301 := "0";
    null;
    r3302 := (r3301);
    r3303 := "0";
    null;
    r3304 := (r3303);
    r3305 := "1";
    null;
    r3306 := (r3305);
    r3307 := "0";
    null;
    r3308 := (r3307);
    r3309 := "0";
    null;
    r3310 := (r3309);
    r3311 := "0";
    null;
    r3312 := (r3311);
    r3313 := "1";
    null;
    r3314 := (r3313);
    r3315 := "1";
    null;
    r3316 := (r3315);
    r3317 := "1";
    null;
    r3318 := (r3317);
    r3319 := "1";
    null;
    r3320 := (r3319);
    r3321 := "1";
    null;
    r3322 := (r3321);
    r3323 := "1";
    null;
    r3324 := (r3323);
    r3325 := "1";
    null;
    r3326 := (r3325);
    r3327 := "0";
    null;
    r3328 := (r3327);
    r3329 := "0";
    null;
    r3330 := (r3329);
    r3331 := "0";
    null;
    r3332 := (r3331);
    r3333 := "0";
    null;
    r3334 := (r3333);
    r3335 := "0";
    null;
    r3336 := (r3335);
    r3337 := "1";
    null;
    r3338 := (r3337);
    r3339 := "0";
    null;
    r3340 := (r3339);
    r3341 := "1";
    null;
    r3342 := (r3341);
    r3343 := "0";
    null;
    r3344 := (r3343);
    r3345 := "1";
    null;
    r3346 := (r3345);
    r3347 := "0";
    null;
    r3348 := (r3347);
    r3349 := "0";
    null;
    r3350 := (r3349);
    r3351 := "1";
    null;
    r3352 := (r3351);
    r3353 := "0";
    null;
    r3354 := (r3353);
    r3355 := "0";
    null;
    r3356 := (r3355);
    r3292 := (r3294 & r3296 & r3298 & r3300 & r3302 & r3304 & r3306 & r3308 & r3310 & r3312 & r3314 & r3316 & r3318 & r3320 & r3322 & r3324 & r3326 & r3328 & r3330 & r3332 & r3334 & r3336 & r3338 & r3340 & r3342 & r3344 & r3346 & r3348 & r3350 & r3352 & r3354 & r3356);
    return r3292;
  end rewire_MetaprogrammingRWw923f82a4_3291;
  function rewire_MetaprogrammingRWw59f111f1_3222 return std_logic_vector
  is
    variable r3287 : std_logic_vector(0 to 0) := (others => '0');
    variable r3286 : std_logic_vector(0 to 0) := (others => '0');
    variable r3285 : std_logic_vector(0 to 0) := (others => '0');
    variable r3284 : std_logic_vector(0 to 0) := (others => '0');
    variable r3283 : std_logic_vector(0 to 0) := (others => '0');
    variable r3282 : std_logic_vector(0 to 0) := (others => '0');
    variable r3281 : std_logic_vector(0 to 0) := (others => '0');
    variable r3280 : std_logic_vector(0 to 0) := (others => '0');
    variable r3279 : std_logic_vector(0 to 0) := (others => '0');
    variable r3278 : std_logic_vector(0 to 0) := (others => '0');
    variable r3277 : std_logic_vector(0 to 0) := (others => '0');
    variable r3276 : std_logic_vector(0 to 0) := (others => '0');
    variable r3275 : std_logic_vector(0 to 0) := (others => '0');
    variable r3274 : std_logic_vector(0 to 0) := (others => '0');
    variable r3273 : std_logic_vector(0 to 0) := (others => '0');
    variable r3272 : std_logic_vector(0 to 0) := (others => '0');
    variable r3271 : std_logic_vector(0 to 0) := (others => '0');
    variable r3270 : std_logic_vector(0 to 0) := (others => '0');
    variable r3269 : std_logic_vector(0 to 0) := (others => '0');
    variable r3268 : std_logic_vector(0 to 0) := (others => '0');
    variable r3267 : std_logic_vector(0 to 0) := (others => '0');
    variable r3266 : std_logic_vector(0 to 0) := (others => '0');
    variable r3265 : std_logic_vector(0 to 0) := (others => '0');
    variable r3264 : std_logic_vector(0 to 0) := (others => '0');
    variable r3263 : std_logic_vector(0 to 0) := (others => '0');
    variable r3262 : std_logic_vector(0 to 0) := (others => '0');
    variable r3261 : std_logic_vector(0 to 0) := (others => '0');
    variable r3260 : std_logic_vector(0 to 0) := (others => '0');
    variable r3259 : std_logic_vector(0 to 0) := (others => '0');
    variable r3258 : std_logic_vector(0 to 0) := (others => '0');
    variable r3257 : std_logic_vector(0 to 0) := (others => '0');
    variable r3256 : std_logic_vector(0 to 0) := (others => '0');
    variable r3255 : std_logic_vector(0 to 0) := (others => '0');
    variable r3254 : std_logic_vector(0 to 0) := (others => '0');
    variable r3253 : std_logic_vector(0 to 0) := (others => '0');
    variable r3252 : std_logic_vector(0 to 0) := (others => '0');
    variable r3251 : std_logic_vector(0 to 0) := (others => '0');
    variable r3250 : std_logic_vector(0 to 0) := (others => '0');
    variable r3249 : std_logic_vector(0 to 0) := (others => '0');
    variable r3248 : std_logic_vector(0 to 0) := (others => '0');
    variable r3247 : std_logic_vector(0 to 0) := (others => '0');
    variable r3246 : std_logic_vector(0 to 0) := (others => '0');
    variable r3245 : std_logic_vector(0 to 0) := (others => '0');
    variable r3244 : std_logic_vector(0 to 0) := (others => '0');
    variable r3243 : std_logic_vector(0 to 0) := (others => '0');
    variable r3242 : std_logic_vector(0 to 0) := (others => '0');
    variable r3241 : std_logic_vector(0 to 0) := (others => '0');
    variable r3240 : std_logic_vector(0 to 0) := (others => '0');
    variable r3239 : std_logic_vector(0 to 0) := (others => '0');
    variable r3238 : std_logic_vector(0 to 0) := (others => '0');
    variable r3237 : std_logic_vector(0 to 0) := (others => '0');
    variable r3236 : std_logic_vector(0 to 0) := (others => '0');
    variable r3235 : std_logic_vector(0 to 0) := (others => '0');
    variable r3234 : std_logic_vector(0 to 0) := (others => '0');
    variable r3233 : std_logic_vector(0 to 0) := (others => '0');
    variable r3232 : std_logic_vector(0 to 0) := (others => '0');
    variable r3231 : std_logic_vector(0 to 0) := (others => '0');
    variable r3230 : std_logic_vector(0 to 0) := (others => '0');
    variable r3229 : std_logic_vector(0 to 0) := (others => '0');
    variable r3228 : std_logic_vector(0 to 0) := (others => '0');
    variable r3227 : std_logic_vector(0 to 0) := (others => '0');
    variable r3226 : std_logic_vector(0 to 0) := (others => '0');
    variable r3225 : std_logic_vector(0 to 0) := (others => '0');
    variable r3224 : std_logic_vector(0 to 0) := (others => '0');
    variable r3223 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r3224 := "0";
    null;
    r3225 := (r3224);
    r3226 := "1";
    null;
    r3227 := (r3226);
    r3228 := "0";
    null;
    r3229 := (r3228);
    r3230 := "1";
    null;
    r3231 := (r3230);
    r3232 := "1";
    null;
    r3233 := (r3232);
    r3234 := "0";
    null;
    r3235 := (r3234);
    r3236 := "0";
    null;
    r3237 := (r3236);
    r3238 := "1";
    null;
    r3239 := (r3238);
    r3240 := "1";
    null;
    r3241 := (r3240);
    r3242 := "1";
    null;
    r3243 := (r3242);
    r3244 := "1";
    null;
    r3245 := (r3244);
    r3246 := "1";
    null;
    r3247 := (r3246);
    r3248 := "0";
    null;
    r3249 := (r3248);
    r3250 := "0";
    null;
    r3251 := (r3250);
    r3252 := "0";
    null;
    r3253 := (r3252);
    r3254 := "1";
    null;
    r3255 := (r3254);
    r3256 := "0";
    null;
    r3257 := (r3256);
    r3258 := "0";
    null;
    r3259 := (r3258);
    r3260 := "0";
    null;
    r3261 := (r3260);
    r3262 := "1";
    null;
    r3263 := (r3262);
    r3264 := "0";
    null;
    r3265 := (r3264);
    r3266 := "0";
    null;
    r3267 := (r3266);
    r3268 := "0";
    null;
    r3269 := (r3268);
    r3270 := "1";
    null;
    r3271 := (r3270);
    r3272 := "1";
    null;
    r3273 := (r3272);
    r3274 := "1";
    null;
    r3275 := (r3274);
    r3276 := "1";
    null;
    r3277 := (r3276);
    r3278 := "1";
    null;
    r3279 := (r3278);
    r3280 := "0";
    null;
    r3281 := (r3280);
    r3282 := "0";
    null;
    r3283 := (r3282);
    r3284 := "0";
    null;
    r3285 := (r3284);
    r3286 := "1";
    null;
    r3287 := (r3286);
    r3223 := (r3225 & r3227 & r3229 & r3231 & r3233 & r3235 & r3237 & r3239 & r3241 & r3243 & r3245 & r3247 & r3249 & r3251 & r3253 & r3255 & r3257 & r3259 & r3261 & r3263 & r3265 & r3267 & r3269 & r3271 & r3273 & r3275 & r3277 & r3279 & r3281 & r3283 & r3285 & r3287);
    return r3223;
  end rewire_MetaprogrammingRWw59f111f1_3222;
  function rewire_MetaprogrammingRWw3956c25b_3153 return std_logic_vector
  is
    variable r3218 : std_logic_vector(0 to 0) := (others => '0');
    variable r3217 : std_logic_vector(0 to 0) := (others => '0');
    variable r3216 : std_logic_vector(0 to 0) := (others => '0');
    variable r3215 : std_logic_vector(0 to 0) := (others => '0');
    variable r3214 : std_logic_vector(0 to 0) := (others => '0');
    variable r3213 : std_logic_vector(0 to 0) := (others => '0');
    variable r3212 : std_logic_vector(0 to 0) := (others => '0');
    variable r3211 : std_logic_vector(0 to 0) := (others => '0');
    variable r3210 : std_logic_vector(0 to 0) := (others => '0');
    variable r3209 : std_logic_vector(0 to 0) := (others => '0');
    variable r3208 : std_logic_vector(0 to 0) := (others => '0');
    variable r3207 : std_logic_vector(0 to 0) := (others => '0');
    variable r3206 : std_logic_vector(0 to 0) := (others => '0');
    variable r3205 : std_logic_vector(0 to 0) := (others => '0');
    variable r3204 : std_logic_vector(0 to 0) := (others => '0');
    variable r3203 : std_logic_vector(0 to 0) := (others => '0');
    variable r3202 : std_logic_vector(0 to 0) := (others => '0');
    variable r3201 : std_logic_vector(0 to 0) := (others => '0');
    variable r3200 : std_logic_vector(0 to 0) := (others => '0');
    variable r3199 : std_logic_vector(0 to 0) := (others => '0');
    variable r3198 : std_logic_vector(0 to 0) := (others => '0');
    variable r3197 : std_logic_vector(0 to 0) := (others => '0');
    variable r3196 : std_logic_vector(0 to 0) := (others => '0');
    variable r3195 : std_logic_vector(0 to 0) := (others => '0');
    variable r3194 : std_logic_vector(0 to 0) := (others => '0');
    variable r3193 : std_logic_vector(0 to 0) := (others => '0');
    variable r3192 : std_logic_vector(0 to 0) := (others => '0');
    variable r3191 : std_logic_vector(0 to 0) := (others => '0');
    variable r3190 : std_logic_vector(0 to 0) := (others => '0');
    variable r3189 : std_logic_vector(0 to 0) := (others => '0');
    variable r3188 : std_logic_vector(0 to 0) := (others => '0');
    variable r3187 : std_logic_vector(0 to 0) := (others => '0');
    variable r3186 : std_logic_vector(0 to 0) := (others => '0');
    variable r3185 : std_logic_vector(0 to 0) := (others => '0');
    variable r3184 : std_logic_vector(0 to 0) := (others => '0');
    variable r3183 : std_logic_vector(0 to 0) := (others => '0');
    variable r3182 : std_logic_vector(0 to 0) := (others => '0');
    variable r3181 : std_logic_vector(0 to 0) := (others => '0');
    variable r3180 : std_logic_vector(0 to 0) := (others => '0');
    variable r3179 : std_logic_vector(0 to 0) := (others => '0');
    variable r3178 : std_logic_vector(0 to 0) := (others => '0');
    variable r3177 : std_logic_vector(0 to 0) := (others => '0');
    variable r3176 : std_logic_vector(0 to 0) := (others => '0');
    variable r3175 : std_logic_vector(0 to 0) := (others => '0');
    variable r3174 : std_logic_vector(0 to 0) := (others => '0');
    variable r3173 : std_logic_vector(0 to 0) := (others => '0');
    variable r3172 : std_logic_vector(0 to 0) := (others => '0');
    variable r3171 : std_logic_vector(0 to 0) := (others => '0');
    variable r3170 : std_logic_vector(0 to 0) := (others => '0');
    variable r3169 : std_logic_vector(0 to 0) := (others => '0');
    variable r3168 : std_logic_vector(0 to 0) := (others => '0');
    variable r3167 : std_logic_vector(0 to 0) := (others => '0');
    variable r3166 : std_logic_vector(0 to 0) := (others => '0');
    variable r3165 : std_logic_vector(0 to 0) := (others => '0');
    variable r3164 : std_logic_vector(0 to 0) := (others => '0');
    variable r3163 : std_logic_vector(0 to 0) := (others => '0');
    variable r3162 : std_logic_vector(0 to 0) := (others => '0');
    variable r3161 : std_logic_vector(0 to 0) := (others => '0');
    variable r3160 : std_logic_vector(0 to 0) := (others => '0');
    variable r3159 : std_logic_vector(0 to 0) := (others => '0');
    variable r3158 : std_logic_vector(0 to 0) := (others => '0');
    variable r3157 : std_logic_vector(0 to 0) := (others => '0');
    variable r3156 : std_logic_vector(0 to 0) := (others => '0');
    variable r3155 : std_logic_vector(0 to 0) := (others => '0');
    variable r3154 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r3155 := "0";
    null;
    r3156 := (r3155);
    r3157 := "0";
    null;
    r3158 := (r3157);
    r3159 := "1";
    null;
    r3160 := (r3159);
    r3161 := "1";
    null;
    r3162 := (r3161);
    r3163 := "1";
    null;
    r3164 := (r3163);
    r3165 := "0";
    null;
    r3166 := (r3165);
    r3167 := "0";
    null;
    r3168 := (r3167);
    r3169 := "1";
    null;
    r3170 := (r3169);
    r3171 := "0";
    null;
    r3172 := (r3171);
    r3173 := "1";
    null;
    r3174 := (r3173);
    r3175 := "0";
    null;
    r3176 := (r3175);
    r3177 := "1";
    null;
    r3178 := (r3177);
    r3179 := "0";
    null;
    r3180 := (r3179);
    r3181 := "1";
    null;
    r3182 := (r3181);
    r3183 := "1";
    null;
    r3184 := (r3183);
    r3185 := "0";
    null;
    r3186 := (r3185);
    r3187 := "1";
    null;
    r3188 := (r3187);
    r3189 := "1";
    null;
    r3190 := (r3189);
    r3191 := "0";
    null;
    r3192 := (r3191);
    r3193 := "0";
    null;
    r3194 := (r3193);
    r3195 := "0";
    null;
    r3196 := (r3195);
    r3197 := "0";
    null;
    r3198 := (r3197);
    r3199 := "1";
    null;
    r3200 := (r3199);
    r3201 := "0";
    null;
    r3202 := (r3201);
    r3203 := "0";
    null;
    r3204 := (r3203);
    r3205 := "1";
    null;
    r3206 := (r3205);
    r3207 := "0";
    null;
    r3208 := (r3207);
    r3209 := "1";
    null;
    r3210 := (r3209);
    r3211 := "1";
    null;
    r3212 := (r3211);
    r3213 := "0";
    null;
    r3214 := (r3213);
    r3215 := "1";
    null;
    r3216 := (r3215);
    r3217 := "1";
    null;
    r3218 := (r3217);
    r3154 := (r3156 & r3158 & r3160 & r3162 & r3164 & r3166 & r3168 & r3170 & r3172 & r3174 & r3176 & r3178 & r3180 & r3182 & r3184 & r3186 & r3188 & r3190 & r3192 & r3194 & r3196 & r3198 & r3200 & r3202 & r3204 & r3206 & r3208 & r3210 & r3212 & r3214 & r3216 & r3218);
    return r3154;
  end rewire_MetaprogrammingRWw3956c25b_3153;
  function rewire_MetaprogrammingRWwe9b5dba5_3084 return std_logic_vector
  is
    variable r3149 : std_logic_vector(0 to 0) := (others => '0');
    variable r3148 : std_logic_vector(0 to 0) := (others => '0');
    variable r3147 : std_logic_vector(0 to 0) := (others => '0');
    variable r3146 : std_logic_vector(0 to 0) := (others => '0');
    variable r3145 : std_logic_vector(0 to 0) := (others => '0');
    variable r3144 : std_logic_vector(0 to 0) := (others => '0');
    variable r3143 : std_logic_vector(0 to 0) := (others => '0');
    variable r3142 : std_logic_vector(0 to 0) := (others => '0');
    variable r3141 : std_logic_vector(0 to 0) := (others => '0');
    variable r3140 : std_logic_vector(0 to 0) := (others => '0');
    variable r3139 : std_logic_vector(0 to 0) := (others => '0');
    variable r3138 : std_logic_vector(0 to 0) := (others => '0');
    variable r3137 : std_logic_vector(0 to 0) := (others => '0');
    variable r3136 : std_logic_vector(0 to 0) := (others => '0');
    variable r3135 : std_logic_vector(0 to 0) := (others => '0');
    variable r3134 : std_logic_vector(0 to 0) := (others => '0');
    variable r3133 : std_logic_vector(0 to 0) := (others => '0');
    variable r3132 : std_logic_vector(0 to 0) := (others => '0');
    variable r3131 : std_logic_vector(0 to 0) := (others => '0');
    variable r3130 : std_logic_vector(0 to 0) := (others => '0');
    variable r3129 : std_logic_vector(0 to 0) := (others => '0');
    variable r3128 : std_logic_vector(0 to 0) := (others => '0');
    variable r3127 : std_logic_vector(0 to 0) := (others => '0');
    variable r3126 : std_logic_vector(0 to 0) := (others => '0');
    variable r3125 : std_logic_vector(0 to 0) := (others => '0');
    variable r3124 : std_logic_vector(0 to 0) := (others => '0');
    variable r3123 : std_logic_vector(0 to 0) := (others => '0');
    variable r3122 : std_logic_vector(0 to 0) := (others => '0');
    variable r3121 : std_logic_vector(0 to 0) := (others => '0');
    variable r3120 : std_logic_vector(0 to 0) := (others => '0');
    variable r3119 : std_logic_vector(0 to 0) := (others => '0');
    variable r3118 : std_logic_vector(0 to 0) := (others => '0');
    variable r3117 : std_logic_vector(0 to 0) := (others => '0');
    variable r3116 : std_logic_vector(0 to 0) := (others => '0');
    variable r3115 : std_logic_vector(0 to 0) := (others => '0');
    variable r3114 : std_logic_vector(0 to 0) := (others => '0');
    variable r3113 : std_logic_vector(0 to 0) := (others => '0');
    variable r3112 : std_logic_vector(0 to 0) := (others => '0');
    variable r3111 : std_logic_vector(0 to 0) := (others => '0');
    variable r3110 : std_logic_vector(0 to 0) := (others => '0');
    variable r3109 : std_logic_vector(0 to 0) := (others => '0');
    variable r3108 : std_logic_vector(0 to 0) := (others => '0');
    variable r3107 : std_logic_vector(0 to 0) := (others => '0');
    variable r3106 : std_logic_vector(0 to 0) := (others => '0');
    variable r3105 : std_logic_vector(0 to 0) := (others => '0');
    variable r3104 : std_logic_vector(0 to 0) := (others => '0');
    variable r3103 : std_logic_vector(0 to 0) := (others => '0');
    variable r3102 : std_logic_vector(0 to 0) := (others => '0');
    variable r3101 : std_logic_vector(0 to 0) := (others => '0');
    variable r3100 : std_logic_vector(0 to 0) := (others => '0');
    variable r3099 : std_logic_vector(0 to 0) := (others => '0');
    variable r3098 : std_logic_vector(0 to 0) := (others => '0');
    variable r3097 : std_logic_vector(0 to 0) := (others => '0');
    variable r3096 : std_logic_vector(0 to 0) := (others => '0');
    variable r3095 : std_logic_vector(0 to 0) := (others => '0');
    variable r3094 : std_logic_vector(0 to 0) := (others => '0');
    variable r3093 : std_logic_vector(0 to 0) := (others => '0');
    variable r3092 : std_logic_vector(0 to 0) := (others => '0');
    variable r3091 : std_logic_vector(0 to 0) := (others => '0');
    variable r3090 : std_logic_vector(0 to 0) := (others => '0');
    variable r3089 : std_logic_vector(0 to 0) := (others => '0');
    variable r3088 : std_logic_vector(0 to 0) := (others => '0');
    variable r3087 : std_logic_vector(0 to 0) := (others => '0');
    variable r3086 : std_logic_vector(0 to 0) := (others => '0');
    variable r3085 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r3086 := "1";
    null;
    r3087 := (r3086);
    r3088 := "1";
    null;
    r3089 := (r3088);
    r3090 := "1";
    null;
    r3091 := (r3090);
    r3092 := "0";
    null;
    r3093 := (r3092);
    r3094 := "1";
    null;
    r3095 := (r3094);
    r3096 := "0";
    null;
    r3097 := (r3096);
    r3098 := "0";
    null;
    r3099 := (r3098);
    r3100 := "1";
    null;
    r3101 := (r3100);
    r3102 := "1";
    null;
    r3103 := (r3102);
    r3104 := "0";
    null;
    r3105 := (r3104);
    r3106 := "1";
    null;
    r3107 := (r3106);
    r3108 := "1";
    null;
    r3109 := (r3108);
    r3110 := "0";
    null;
    r3111 := (r3110);
    r3112 := "1";
    null;
    r3113 := (r3112);
    r3114 := "0";
    null;
    r3115 := (r3114);
    r3116 := "1";
    null;
    r3117 := (r3116);
    r3118 := "1";
    null;
    r3119 := (r3118);
    r3120 := "1";
    null;
    r3121 := (r3120);
    r3122 := "0";
    null;
    r3123 := (r3122);
    r3124 := "1";
    null;
    r3125 := (r3124);
    r3126 := "1";
    null;
    r3127 := (r3126);
    r3128 := "0";
    null;
    r3129 := (r3128);
    r3130 := "1";
    null;
    r3131 := (r3130);
    r3132 := "1";
    null;
    r3133 := (r3132);
    r3134 := "1";
    null;
    r3135 := (r3134);
    r3136 := "0";
    null;
    r3137 := (r3136);
    r3138 := "1";
    null;
    r3139 := (r3138);
    r3140 := "0";
    null;
    r3141 := (r3140);
    r3142 := "0";
    null;
    r3143 := (r3142);
    r3144 := "1";
    null;
    r3145 := (r3144);
    r3146 := "0";
    null;
    r3147 := (r3146);
    r3148 := "1";
    null;
    r3149 := (r3148);
    r3085 := (r3087 & r3089 & r3091 & r3093 & r3095 & r3097 & r3099 & r3101 & r3103 & r3105 & r3107 & r3109 & r3111 & r3113 & r3115 & r3117 & r3119 & r3121 & r3123 & r3125 & r3127 & r3129 & r3131 & r3133 & r3135 & r3137 & r3139 & r3141 & r3143 & r3145 & r3147 & r3149);
    return r3085;
  end rewire_MetaprogrammingRWwe9b5dba5_3084;
  function rewire_MetaprogrammingRWwb5c0fbcf_3015 return std_logic_vector
  is
    variable r3080 : std_logic_vector(0 to 0) := (others => '0');
    variable r3079 : std_logic_vector(0 to 0) := (others => '0');
    variable r3078 : std_logic_vector(0 to 0) := (others => '0');
    variable r3077 : std_logic_vector(0 to 0) := (others => '0');
    variable r3076 : std_logic_vector(0 to 0) := (others => '0');
    variable r3075 : std_logic_vector(0 to 0) := (others => '0');
    variable r3074 : std_logic_vector(0 to 0) := (others => '0');
    variable r3073 : std_logic_vector(0 to 0) := (others => '0');
    variable r3072 : std_logic_vector(0 to 0) := (others => '0');
    variable r3071 : std_logic_vector(0 to 0) := (others => '0');
    variable r3070 : std_logic_vector(0 to 0) := (others => '0');
    variable r3069 : std_logic_vector(0 to 0) := (others => '0');
    variable r3068 : std_logic_vector(0 to 0) := (others => '0');
    variable r3067 : std_logic_vector(0 to 0) := (others => '0');
    variable r3066 : std_logic_vector(0 to 0) := (others => '0');
    variable r3065 : std_logic_vector(0 to 0) := (others => '0');
    variable r3064 : std_logic_vector(0 to 0) := (others => '0');
    variable r3063 : std_logic_vector(0 to 0) := (others => '0');
    variable r3062 : std_logic_vector(0 to 0) := (others => '0');
    variable r3061 : std_logic_vector(0 to 0) := (others => '0');
    variable r3060 : std_logic_vector(0 to 0) := (others => '0');
    variable r3059 : std_logic_vector(0 to 0) := (others => '0');
    variable r3058 : std_logic_vector(0 to 0) := (others => '0');
    variable r3057 : std_logic_vector(0 to 0) := (others => '0');
    variable r3056 : std_logic_vector(0 to 0) := (others => '0');
    variable r3055 : std_logic_vector(0 to 0) := (others => '0');
    variable r3054 : std_logic_vector(0 to 0) := (others => '0');
    variable r3053 : std_logic_vector(0 to 0) := (others => '0');
    variable r3052 : std_logic_vector(0 to 0) := (others => '0');
    variable r3051 : std_logic_vector(0 to 0) := (others => '0');
    variable r3050 : std_logic_vector(0 to 0) := (others => '0');
    variable r3049 : std_logic_vector(0 to 0) := (others => '0');
    variable r3048 : std_logic_vector(0 to 0) := (others => '0');
    variable r3047 : std_logic_vector(0 to 0) := (others => '0');
    variable r3046 : std_logic_vector(0 to 0) := (others => '0');
    variable r3045 : std_logic_vector(0 to 0) := (others => '0');
    variable r3044 : std_logic_vector(0 to 0) := (others => '0');
    variable r3043 : std_logic_vector(0 to 0) := (others => '0');
    variable r3042 : std_logic_vector(0 to 0) := (others => '0');
    variable r3041 : std_logic_vector(0 to 0) := (others => '0');
    variable r3040 : std_logic_vector(0 to 0) := (others => '0');
    variable r3039 : std_logic_vector(0 to 0) := (others => '0');
    variable r3038 : std_logic_vector(0 to 0) := (others => '0');
    variable r3037 : std_logic_vector(0 to 0) := (others => '0');
    variable r3036 : std_logic_vector(0 to 0) := (others => '0');
    variable r3035 : std_logic_vector(0 to 0) := (others => '0');
    variable r3034 : std_logic_vector(0 to 0) := (others => '0');
    variable r3033 : std_logic_vector(0 to 0) := (others => '0');
    variable r3032 : std_logic_vector(0 to 0) := (others => '0');
    variable r3031 : std_logic_vector(0 to 0) := (others => '0');
    variable r3030 : std_logic_vector(0 to 0) := (others => '0');
    variable r3029 : std_logic_vector(0 to 0) := (others => '0');
    variable r3028 : std_logic_vector(0 to 0) := (others => '0');
    variable r3027 : std_logic_vector(0 to 0) := (others => '0');
    variable r3026 : std_logic_vector(0 to 0) := (others => '0');
    variable r3025 : std_logic_vector(0 to 0) := (others => '0');
    variable r3024 : std_logic_vector(0 to 0) := (others => '0');
    variable r3023 : std_logic_vector(0 to 0) := (others => '0');
    variable r3022 : std_logic_vector(0 to 0) := (others => '0');
    variable r3021 : std_logic_vector(0 to 0) := (others => '0');
    variable r3020 : std_logic_vector(0 to 0) := (others => '0');
    variable r3019 : std_logic_vector(0 to 0) := (others => '0');
    variable r3018 : std_logic_vector(0 to 0) := (others => '0');
    variable r3017 : std_logic_vector(0 to 0) := (others => '0');
    variable r3016 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r3017 := "1";
    null;
    r3018 := (r3017);
    r3019 := "0";
    null;
    r3020 := (r3019);
    r3021 := "1";
    null;
    r3022 := (r3021);
    r3023 := "1";
    null;
    r3024 := (r3023);
    r3025 := "0";
    null;
    r3026 := (r3025);
    r3027 := "1";
    null;
    r3028 := (r3027);
    r3029 := "0";
    null;
    r3030 := (r3029);
    r3031 := "1";
    null;
    r3032 := (r3031);
    r3033 := "1";
    null;
    r3034 := (r3033);
    r3035 := "1";
    null;
    r3036 := (r3035);
    r3037 := "0";
    null;
    r3038 := (r3037);
    r3039 := "0";
    null;
    r3040 := (r3039);
    r3041 := "0";
    null;
    r3042 := (r3041);
    r3043 := "0";
    null;
    r3044 := (r3043);
    r3045 := "0";
    null;
    r3046 := (r3045);
    r3047 := "0";
    null;
    r3048 := (r3047);
    r3049 := "1";
    null;
    r3050 := (r3049);
    r3051 := "1";
    null;
    r3052 := (r3051);
    r3053 := "1";
    null;
    r3054 := (r3053);
    r3055 := "1";
    null;
    r3056 := (r3055);
    r3057 := "1";
    null;
    r3058 := (r3057);
    r3059 := "0";
    null;
    r3060 := (r3059);
    r3061 := "1";
    null;
    r3062 := (r3061);
    r3063 := "1";
    null;
    r3064 := (r3063);
    r3065 := "1";
    null;
    r3066 := (r3065);
    r3067 := "1";
    null;
    r3068 := (r3067);
    r3069 := "0";
    null;
    r3070 := (r3069);
    r3071 := "0";
    null;
    r3072 := (r3071);
    r3073 := "1";
    null;
    r3074 := (r3073);
    r3075 := "1";
    null;
    r3076 := (r3075);
    r3077 := "1";
    null;
    r3078 := (r3077);
    r3079 := "1";
    null;
    r3080 := (r3079);
    r3016 := (r3018 & r3020 & r3022 & r3024 & r3026 & r3028 & r3030 & r3032 & r3034 & r3036 & r3038 & r3040 & r3042 & r3044 & r3046 & r3048 & r3050 & r3052 & r3054 & r3056 & r3058 & r3060 & r3062 & r3064 & r3066 & r3068 & r3070 & r3072 & r3074 & r3076 & r3078 & r3080);
    return r3016;
  end rewire_MetaprogrammingRWwb5c0fbcf_3015;
  function rewire_MetaprogrammingRWw71374491_2946 return std_logic_vector
  is
    variable r3011 : std_logic_vector(0 to 0) := (others => '0');
    variable r3010 : std_logic_vector(0 to 0) := (others => '0');
    variable r3009 : std_logic_vector(0 to 0) := (others => '0');
    variable r3008 : std_logic_vector(0 to 0) := (others => '0');
    variable r3007 : std_logic_vector(0 to 0) := (others => '0');
    variable r3006 : std_logic_vector(0 to 0) := (others => '0');
    variable r3005 : std_logic_vector(0 to 0) := (others => '0');
    variable r3004 : std_logic_vector(0 to 0) := (others => '0');
    variable r3003 : std_logic_vector(0 to 0) := (others => '0');
    variable r3002 : std_logic_vector(0 to 0) := (others => '0');
    variable r3001 : std_logic_vector(0 to 0) := (others => '0');
    variable r3000 : std_logic_vector(0 to 0) := (others => '0');
    variable r2999 : std_logic_vector(0 to 0) := (others => '0');
    variable r2998 : std_logic_vector(0 to 0) := (others => '0');
    variable r2997 : std_logic_vector(0 to 0) := (others => '0');
    variable r2996 : std_logic_vector(0 to 0) := (others => '0');
    variable r2995 : std_logic_vector(0 to 0) := (others => '0');
    variable r2994 : std_logic_vector(0 to 0) := (others => '0');
    variable r2993 : std_logic_vector(0 to 0) := (others => '0');
    variable r2992 : std_logic_vector(0 to 0) := (others => '0');
    variable r2991 : std_logic_vector(0 to 0) := (others => '0');
    variable r2990 : std_logic_vector(0 to 0) := (others => '0');
    variable r2989 : std_logic_vector(0 to 0) := (others => '0');
    variable r2988 : std_logic_vector(0 to 0) := (others => '0');
    variable r2987 : std_logic_vector(0 to 0) := (others => '0');
    variable r2986 : std_logic_vector(0 to 0) := (others => '0');
    variable r2985 : std_logic_vector(0 to 0) := (others => '0');
    variable r2984 : std_logic_vector(0 to 0) := (others => '0');
    variable r2983 : std_logic_vector(0 to 0) := (others => '0');
    variable r2982 : std_logic_vector(0 to 0) := (others => '0');
    variable r2981 : std_logic_vector(0 to 0) := (others => '0');
    variable r2980 : std_logic_vector(0 to 0) := (others => '0');
    variable r2979 : std_logic_vector(0 to 0) := (others => '0');
    variable r2978 : std_logic_vector(0 to 0) := (others => '0');
    variable r2977 : std_logic_vector(0 to 0) := (others => '0');
    variable r2976 : std_logic_vector(0 to 0) := (others => '0');
    variable r2975 : std_logic_vector(0 to 0) := (others => '0');
    variable r2974 : std_logic_vector(0 to 0) := (others => '0');
    variable r2973 : std_logic_vector(0 to 0) := (others => '0');
    variable r2972 : std_logic_vector(0 to 0) := (others => '0');
    variable r2971 : std_logic_vector(0 to 0) := (others => '0');
    variable r2970 : std_logic_vector(0 to 0) := (others => '0');
    variable r2969 : std_logic_vector(0 to 0) := (others => '0');
    variable r2968 : std_logic_vector(0 to 0) := (others => '0');
    variable r2967 : std_logic_vector(0 to 0) := (others => '0');
    variable r2966 : std_logic_vector(0 to 0) := (others => '0');
    variable r2965 : std_logic_vector(0 to 0) := (others => '0');
    variable r2964 : std_logic_vector(0 to 0) := (others => '0');
    variable r2963 : std_logic_vector(0 to 0) := (others => '0');
    variable r2962 : std_logic_vector(0 to 0) := (others => '0');
    variable r2961 : std_logic_vector(0 to 0) := (others => '0');
    variable r2960 : std_logic_vector(0 to 0) := (others => '0');
    variable r2959 : std_logic_vector(0 to 0) := (others => '0');
    variable r2958 : std_logic_vector(0 to 0) := (others => '0');
    variable r2957 : std_logic_vector(0 to 0) := (others => '0');
    variable r2956 : std_logic_vector(0 to 0) := (others => '0');
    variable r2955 : std_logic_vector(0 to 0) := (others => '0');
    variable r2954 : std_logic_vector(0 to 0) := (others => '0');
    variable r2953 : std_logic_vector(0 to 0) := (others => '0');
    variable r2952 : std_logic_vector(0 to 0) := (others => '0');
    variable r2951 : std_logic_vector(0 to 0) := (others => '0');
    variable r2950 : std_logic_vector(0 to 0) := (others => '0');
    variable r2949 : std_logic_vector(0 to 0) := (others => '0');
    variable r2948 : std_logic_vector(0 to 0) := (others => '0');
    variable r2947 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r2948 := "0";
    null;
    r2949 := (r2948);
    r2950 := "1";
    null;
    r2951 := (r2950);
    r2952 := "1";
    null;
    r2953 := (r2952);
    r2954 := "1";
    null;
    r2955 := (r2954);
    r2956 := "0";
    null;
    r2957 := (r2956);
    r2958 := "0";
    null;
    r2959 := (r2958);
    r2960 := "0";
    null;
    r2961 := (r2960);
    r2962 := "1";
    null;
    r2963 := (r2962);
    r2964 := "0";
    null;
    r2965 := (r2964);
    r2966 := "0";
    null;
    r2967 := (r2966);
    r2968 := "1";
    null;
    r2969 := (r2968);
    r2970 := "1";
    null;
    r2971 := (r2970);
    r2972 := "0";
    null;
    r2973 := (r2972);
    r2974 := "1";
    null;
    r2975 := (r2974);
    r2976 := "1";
    null;
    r2977 := (r2976);
    r2978 := "1";
    null;
    r2979 := (r2978);
    r2980 := "0";
    null;
    r2981 := (r2980);
    r2982 := "1";
    null;
    r2983 := (r2982);
    r2984 := "0";
    null;
    r2985 := (r2984);
    r2986 := "0";
    null;
    r2987 := (r2986);
    r2988 := "0";
    null;
    r2989 := (r2988);
    r2990 := "1";
    null;
    r2991 := (r2990);
    r2992 := "0";
    null;
    r2993 := (r2992);
    r2994 := "0";
    null;
    r2995 := (r2994);
    r2996 := "1";
    null;
    r2997 := (r2996);
    r2998 := "0";
    null;
    r2999 := (r2998);
    r3000 := "0";
    null;
    r3001 := (r3000);
    r3002 := "1";
    null;
    r3003 := (r3002);
    r3004 := "0";
    null;
    r3005 := (r3004);
    r3006 := "0";
    null;
    r3007 := (r3006);
    r3008 := "0";
    null;
    r3009 := (r3008);
    r3010 := "1";
    null;
    r3011 := (r3010);
    r2947 := (r2949 & r2951 & r2953 & r2955 & r2957 & r2959 & r2961 & r2963 & r2965 & r2967 & r2969 & r2971 & r2973 & r2975 & r2977 & r2979 & r2981 & r2983 & r2985 & r2987 & r2989 & r2991 & r2993 & r2995 & r2997 & r2999 & r3001 & r3003 & r3005 & r3007 & r3009 & r3011);
    return r2947;
  end rewire_MetaprogrammingRWw71374491_2946;
  function rewire_MetaprogrammingRWw428a2f98_2877 return std_logic_vector
  is
    variable r2942 : std_logic_vector(0 to 0) := (others => '0');
    variable r2941 : std_logic_vector(0 to 0) := (others => '0');
    variable r2940 : std_logic_vector(0 to 0) := (others => '0');
    variable r2939 : std_logic_vector(0 to 0) := (others => '0');
    variable r2938 : std_logic_vector(0 to 0) := (others => '0');
    variable r2937 : std_logic_vector(0 to 0) := (others => '0');
    variable r2936 : std_logic_vector(0 to 0) := (others => '0');
    variable r2935 : std_logic_vector(0 to 0) := (others => '0');
    variable r2934 : std_logic_vector(0 to 0) := (others => '0');
    variable r2933 : std_logic_vector(0 to 0) := (others => '0');
    variable r2932 : std_logic_vector(0 to 0) := (others => '0');
    variable r2931 : std_logic_vector(0 to 0) := (others => '0');
    variable r2930 : std_logic_vector(0 to 0) := (others => '0');
    variable r2929 : std_logic_vector(0 to 0) := (others => '0');
    variable r2928 : std_logic_vector(0 to 0) := (others => '0');
    variable r2927 : std_logic_vector(0 to 0) := (others => '0');
    variable r2926 : std_logic_vector(0 to 0) := (others => '0');
    variable r2925 : std_logic_vector(0 to 0) := (others => '0');
    variable r2924 : std_logic_vector(0 to 0) := (others => '0');
    variable r2923 : std_logic_vector(0 to 0) := (others => '0');
    variable r2922 : std_logic_vector(0 to 0) := (others => '0');
    variable r2921 : std_logic_vector(0 to 0) := (others => '0');
    variable r2920 : std_logic_vector(0 to 0) := (others => '0');
    variable r2919 : std_logic_vector(0 to 0) := (others => '0');
    variable r2918 : std_logic_vector(0 to 0) := (others => '0');
    variable r2917 : std_logic_vector(0 to 0) := (others => '0');
    variable r2916 : std_logic_vector(0 to 0) := (others => '0');
    variable r2915 : std_logic_vector(0 to 0) := (others => '0');
    variable r2914 : std_logic_vector(0 to 0) := (others => '0');
    variable r2913 : std_logic_vector(0 to 0) := (others => '0');
    variable r2912 : std_logic_vector(0 to 0) := (others => '0');
    variable r2911 : std_logic_vector(0 to 0) := (others => '0');
    variable r2910 : std_logic_vector(0 to 0) := (others => '0');
    variable r2909 : std_logic_vector(0 to 0) := (others => '0');
    variable r2908 : std_logic_vector(0 to 0) := (others => '0');
    variable r2907 : std_logic_vector(0 to 0) := (others => '0');
    variable r2906 : std_logic_vector(0 to 0) := (others => '0');
    variable r2905 : std_logic_vector(0 to 0) := (others => '0');
    variable r2904 : std_logic_vector(0 to 0) := (others => '0');
    variable r2903 : std_logic_vector(0 to 0) := (others => '0');
    variable r2902 : std_logic_vector(0 to 0) := (others => '0');
    variable r2901 : std_logic_vector(0 to 0) := (others => '0');
    variable r2900 : std_logic_vector(0 to 0) := (others => '0');
    variable r2899 : std_logic_vector(0 to 0) := (others => '0');
    variable r2898 : std_logic_vector(0 to 0) := (others => '0');
    variable r2897 : std_logic_vector(0 to 0) := (others => '0');
    variable r2896 : std_logic_vector(0 to 0) := (others => '0');
    variable r2895 : std_logic_vector(0 to 0) := (others => '0');
    variable r2894 : std_logic_vector(0 to 0) := (others => '0');
    variable r2893 : std_logic_vector(0 to 0) := (others => '0');
    variable r2892 : std_logic_vector(0 to 0) := (others => '0');
    variable r2891 : std_logic_vector(0 to 0) := (others => '0');
    variable r2890 : std_logic_vector(0 to 0) := (others => '0');
    variable r2889 : std_logic_vector(0 to 0) := (others => '0');
    variable r2888 : std_logic_vector(0 to 0) := (others => '0');
    variable r2887 : std_logic_vector(0 to 0) := (others => '0');
    variable r2886 : std_logic_vector(0 to 0) := (others => '0');
    variable r2885 : std_logic_vector(0 to 0) := (others => '0');
    variable r2884 : std_logic_vector(0 to 0) := (others => '0');
    variable r2883 : std_logic_vector(0 to 0) := (others => '0');
    variable r2882 : std_logic_vector(0 to 0) := (others => '0');
    variable r2881 : std_logic_vector(0 to 0) := (others => '0');
    variable r2880 : std_logic_vector(0 to 0) := (others => '0');
    variable r2879 : std_logic_vector(0 to 0) := (others => '0');
    variable r2878 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r2879 := "0";
    null;
    r2880 := (r2879);
    r2881 := "1";
    null;
    r2882 := (r2881);
    r2883 := "0";
    null;
    r2884 := (r2883);
    r2885 := "0";
    null;
    r2886 := (r2885);
    r2887 := "0";
    null;
    r2888 := (r2887);
    r2889 := "0";
    null;
    r2890 := (r2889);
    r2891 := "1";
    null;
    r2892 := (r2891);
    r2893 := "0";
    null;
    r2894 := (r2893);
    r2895 := "1";
    null;
    r2896 := (r2895);
    r2897 := "0";
    null;
    r2898 := (r2897);
    r2899 := "0";
    null;
    r2900 := (r2899);
    r2901 := "0";
    null;
    r2902 := (r2901);
    r2903 := "1";
    null;
    r2904 := (r2903);
    r2905 := "0";
    null;
    r2906 := (r2905);
    r2907 := "1";
    null;
    r2908 := (r2907);
    r2909 := "0";
    null;
    r2910 := (r2909);
    r2911 := "0";
    null;
    r2912 := (r2911);
    r2913 := "0";
    null;
    r2914 := (r2913);
    r2915 := "1";
    null;
    r2916 := (r2915);
    r2917 := "0";
    null;
    r2918 := (r2917);
    r2919 := "1";
    null;
    r2920 := (r2919);
    r2921 := "1";
    null;
    r2922 := (r2921);
    r2923 := "1";
    null;
    r2924 := (r2923);
    r2925 := "1";
    null;
    r2926 := (r2925);
    r2927 := "1";
    null;
    r2928 := (r2927);
    r2929 := "0";
    null;
    r2930 := (r2929);
    r2931 := "0";
    null;
    r2932 := (r2931);
    r2933 := "1";
    null;
    r2934 := (r2933);
    r2935 := "1";
    null;
    r2936 := (r2935);
    r2937 := "0";
    null;
    r2938 := (r2937);
    r2939 := "0";
    null;
    r2940 := (r2939);
    r2941 := "0";
    null;
    r2942 := (r2941);
    r2878 := (r2880 & r2882 & r2884 & r2886 & r2888 & r2890 & r2892 & r2894 & r2896 & r2898 & r2900 & r2902 & r2904 & r2906 & r2908 & r2910 & r2912 & r2914 & r2916 & r2918 & r2920 & r2922 & r2924 & r2926 & r2928 & r2930 & r2932 & r2934 & r2936 & r2938 & r2940 & r2942);
    return r2878;
  end rewire_MetaprogrammingRWw428a2f98_2877;
  function rewire_Mainstep256_2373(r2374 : std_logic_vector ; r2375 : std_logic_vector ; r2376 : std_logic_vector) return std_logic_vector
  is
    variable r2872 : std_logic_vector(0 to 31) := (others => '0');
    variable r2871 : std_logic_vector(0 to 31) := (others => '0');
    variable r2870 : std_logic_vector(0 to 31) := (others => '0');
    variable r2869 : std_logic_vector(0 to 31) := (others => '0');
    variable r2868 : std_logic_vector(0 to 31) := (others => '0');
    variable r2867 : std_logic_vector(0 to 31) := (others => '0');
    variable r2866 : std_logic_vector(0 to 31) := (others => '0');
    variable r2865 : std_logic_vector(0 to 31) := (others => '0');
    variable r2864 : std_logic_vector(0 to 31) := (others => '0');
    variable r2863 : std_logic_vector(0 to 31) := (others => '0');
    variable r2857 : std_logic_vector(0 to 31) := (others => '0');
    variable r2856 : std_logic_vector(0 to 31) := (others => '0');
    variable r2855 : std_logic_vector(0 to 31) := (others => '0');
    variable r2853 : std_logic_vector(0 to 31) := (others => '0');
    variable r2637 : std_logic_vector(0 to 31) := (others => '0');
    variable r2635 : std_logic_vector(0 to 31) := (others => '0');
    variable r2634 : std_logic_vector(0 to 31) := (others => '0');
    variable r2633 : std_logic_vector(0 to 31) := (others => '0');
    variable r2632 : std_logic_vector(0 to 31) := (others => '0');
    variable r2631 : std_logic_vector(0 to 31) := (others => '0');
    variable r2626 : std_logic_vector(0 to 31) := (others => '0');
    variable r2625 : std_logic_vector(0 to 31) := (others => '0');
    variable r2624 : std_logic_vector(0 to 31) := (others => '0');
    variable r2622 : std_logic_vector(0 to 31) := (others => '0');
    variable r2406 : std_logic_vector(0 to 31) := (others => '0');
    variable r2404 : std_logic_vector(0 to 255) := (others => '0');
    variable b2403 : boolean := false;
    variable b2402 : boolean := false;
    variable b2401 : boolean := false;
    variable b2400 : boolean := false;
    variable b2399 : boolean := false;
    variable b2398 : boolean := false;
    variable b2397 : boolean := false;
    variable b2396 : boolean := false;
    variable b2395 : boolean := false;
    variable b2394 : boolean := false;
    variable r2393 : std_logic_vector(0 to 31) := (others => '0');
    variable r2392 : std_logic_vector(0 to 31) := (others => '0');
    variable r2391 : std_logic_vector(0 to 31) := (others => '0');
    variable r2390 : std_logic_vector(0 to 31) := (others => '0');
    variable r2389 : std_logic_vector(0 to 31) := (others => '0');
    variable r2388 : std_logic_vector(0 to 31) := (others => '0');
    variable r2387 : std_logic_vector(0 to 31) := (others => '0');
    variable r2386 : std_logic_vector(0 to 31) := (others => '0');
    variable b2385 : boolean := false;
    variable b2384 : boolean := false;
    variable b2383 : boolean := false;
    variable r2382 : std_logic_vector(0 to 255) := (others => '0');
    variable r2381 : std_logic_vector(0 to 31) := (others => '0');
    variable r2380 : std_logic_vector(0 to 31) := (others => '0');
    variable b2379 : boolean := false;
    variable r2378 : std_logic_vector(0 to 255) := (others => '0');
    variable r2377 : std_logic_vector(0 to 319) := (others => '0');
  begin
    null;
    null;
    null;
    null;
    null;
    r2377 := (r2374 & r2375 & r2376);
    b2379 := true;
    r2380 := r2377(0 to 31);
    r2381 := r2377(32 to 63);
    r2382 := r2377(64 to 319);
    b2383 := true;
    b2384 := true;
    b2385 := true;
    r2386 := r2382(0 to 31);
    r2387 := r2382(32 to 63);
    r2388 := r2382(64 to 95);
    r2389 := r2382(96 to 127);
    r2390 := r2382(128 to 159);
    r2391 := r2382(160 to 191);
    r2392 := r2382(192 to 223);
    r2393 := r2382(224 to 255);
    b2394 := true;
    b2395 := true;
    b2396 := true;
    b2397 := true;
    b2398 := true;
    b2399 := true;
    b2400 := true;
    b2401 := true;
    b2402 := (b2385 AND (b2394 AND (b2395 AND (b2396 AND (b2397 AND (b2398 AND (b2399 AND (b2400 AND b2401))))))));
    b2403 := (b2379 AND (b2383 AND (b2384 AND b2402)));
    null;
    null;
    null;
    null;
    r2622 := rewire_Mainbigsigma1_2405(r2390);
    null;
    null;
    null;
    r2631 := rewire_Mainch_2623(r2390,r2391,r2392);
    r2632 := w32Plus(r2622,r2631);
    null;
    null;
    r2633 := w32Plus(r2380,r2381);
    r2634 := w32Plus(r2632,r2633);
    r2635 := w32Plus(r2393,r2634);
    null;
    r2853 := rewire_Mainbigsigma0_2636(r2386);
    null;
    null;
    null;
    r2863 := rewire_Mainmaj_2854(r2386,r2387,r2388);
    r2864 := w32Plus(r2853,r2863);
    r2865 := w32Plus(r2635,r2864);
    null;
    null;
    null;
    null;
    null;
    null;
    r2866 := rewire_Mainbigsigma1_2405(r2390);
    null;
    null;
    null;
    r2867 := rewire_Mainch_2623(r2390,r2391,r2392);
    r2868 := w32Plus(r2866,r2867);
    null;
    null;
    r2869 := w32Plus(r2380,r2381);
    r2870 := w32Plus(r2868,r2869);
    r2871 := w32Plus(r2393,r2870);
    r2872 := w32Plus(r2389,r2871);
    null;
    null;
    null;
    r2404 := (r2865 & r2386 & r2387 & r2388 & r2872 & r2390 & r2391 & r2392);
    r2378 := r2404;
    return r2378;
  end rewire_Mainstep256_2373;
  function rewire_Mainmaj_2854(r2855 : std_logic_vector ; r2856 : std_logic_vector ; r2857 : std_logic_vector) return std_logic_vector
  is
    variable r2862 : std_logic_vector(0 to 31) := (others => '0');
    variable r2861 : std_logic_vector(0 to 31) := (others => '0');
    variable r2860 : std_logic_vector(0 to 31) := (others => '0');
    variable r2859 : std_logic_vector(0 to 31) := (others => '0');
    variable r2858 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r2858 := w32And(r2855,r2856);
    null;
    null;
    r2859 := w32And(r2855,r2857);
    r2860 := w32Xor(r2858,r2859);
    null;
    null;
    r2861 := w32And(r2856,r2857);
    r2862 := w32Xor(r2860,r2861);
    return r2862;
  end rewire_Mainmaj_2854;
  function rewire_Mainbigsigma0_2636(r2637 : std_logic_vector) return std_logic_vector
  is
    variable r2852 : std_logic_vector(0 to 31) := (others => '0');
    variable r2851 : std_logic_vector(0 to 31) := (others => '0');
    variable r2782 : std_logic_vector(0 to 31) := (others => '0');
    variable r2780 : std_logic_vector(0 to 31) := (others => '0');
    variable r2779 : std_logic_vector(0 to 31) := (others => '0');
    variable r2710 : std_logic_vector(0 to 31) := (others => '0');
    variable r2708 : std_logic_vector(0 to 31) := (others => '0');
    variable r2639 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    r2708 := rewire_RWPreluderotateR2_2638(r2637);
    null;
    r2779 := rewire_RWPreluderotateR13_2709(r2637);
    r2780 := w32Xor(r2708,r2779);
    null;
    r2851 := rewire_RWPreluderotateR22_2781(r2637);
    r2852 := w32Xor(r2780,r2851);
    return r2852;
  end rewire_Mainbigsigma0_2636;
  function rewire_RWPreluderotateR22_2781(r2782 : std_logic_vector) return std_logic_vector
  is
    variable r2850 : std_logic_vector(0 to 31) := (others => '0');
    variable b2849 : boolean := false;
    variable b2848 : boolean := false;
    variable b2847 : boolean := false;
    variable b2846 : boolean := false;
    variable b2845 : boolean := false;
    variable b2844 : boolean := false;
    variable b2843 : boolean := false;
    variable b2842 : boolean := false;
    variable b2841 : boolean := false;
    variable b2840 : boolean := false;
    variable b2839 : boolean := false;
    variable b2838 : boolean := false;
    variable b2837 : boolean := false;
    variable b2836 : boolean := false;
    variable b2835 : boolean := false;
    variable b2834 : boolean := false;
    variable b2833 : boolean := false;
    variable b2832 : boolean := false;
    variable b2831 : boolean := false;
    variable b2830 : boolean := false;
    variable b2829 : boolean := false;
    variable b2828 : boolean := false;
    variable b2827 : boolean := false;
    variable b2826 : boolean := false;
    variable b2825 : boolean := false;
    variable b2824 : boolean := false;
    variable b2823 : boolean := false;
    variable b2822 : boolean := false;
    variable b2821 : boolean := false;
    variable b2820 : boolean := false;
    variable b2819 : boolean := false;
    variable b2818 : boolean := false;
    variable b2817 : boolean := false;
    variable r2816 : std_logic_vector(0 to 0) := (others => '0');
    variable r2815 : std_logic_vector(0 to 0) := (others => '0');
    variable r2814 : std_logic_vector(0 to 0) := (others => '0');
    variable r2813 : std_logic_vector(0 to 0) := (others => '0');
    variable r2812 : std_logic_vector(0 to 0) := (others => '0');
    variable r2811 : std_logic_vector(0 to 0) := (others => '0');
    variable r2810 : std_logic_vector(0 to 0) := (others => '0');
    variable r2809 : std_logic_vector(0 to 0) := (others => '0');
    variable r2808 : std_logic_vector(0 to 0) := (others => '0');
    variable r2807 : std_logic_vector(0 to 0) := (others => '0');
    variable r2806 : std_logic_vector(0 to 0) := (others => '0');
    variable r2805 : std_logic_vector(0 to 0) := (others => '0');
    variable r2804 : std_logic_vector(0 to 0) := (others => '0');
    variable r2803 : std_logic_vector(0 to 0) := (others => '0');
    variable r2802 : std_logic_vector(0 to 0) := (others => '0');
    variable r2801 : std_logic_vector(0 to 0) := (others => '0');
    variable r2800 : std_logic_vector(0 to 0) := (others => '0');
    variable r2799 : std_logic_vector(0 to 0) := (others => '0');
    variable r2798 : std_logic_vector(0 to 0) := (others => '0');
    variable r2797 : std_logic_vector(0 to 0) := (others => '0');
    variable r2796 : std_logic_vector(0 to 0) := (others => '0');
    variable r2795 : std_logic_vector(0 to 0) := (others => '0');
    variable r2794 : std_logic_vector(0 to 0) := (others => '0');
    variable r2793 : std_logic_vector(0 to 0) := (others => '0');
    variable r2792 : std_logic_vector(0 to 0) := (others => '0');
    variable r2791 : std_logic_vector(0 to 0) := (others => '0');
    variable r2790 : std_logic_vector(0 to 0) := (others => '0');
    variable r2789 : std_logic_vector(0 to 0) := (others => '0');
    variable r2788 : std_logic_vector(0 to 0) := (others => '0');
    variable r2787 : std_logic_vector(0 to 0) := (others => '0');
    variable r2786 : std_logic_vector(0 to 0) := (others => '0');
    variable r2785 : std_logic_vector(0 to 0) := (others => '0');
    variable b2784 : boolean := false;
    variable r2783 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    b2784 := true;
    r2785 := r2782(0 to 0);
    r2786 := r2782(1 to 1);
    r2787 := r2782(2 to 2);
    r2788 := r2782(3 to 3);
    r2789 := r2782(4 to 4);
    r2790 := r2782(5 to 5);
    r2791 := r2782(6 to 6);
    r2792 := r2782(7 to 7);
    r2793 := r2782(8 to 8);
    r2794 := r2782(9 to 9);
    r2795 := r2782(10 to 10);
    r2796 := r2782(11 to 11);
    r2797 := r2782(12 to 12);
    r2798 := r2782(13 to 13);
    r2799 := r2782(14 to 14);
    r2800 := r2782(15 to 15);
    r2801 := r2782(16 to 16);
    r2802 := r2782(17 to 17);
    r2803 := r2782(18 to 18);
    r2804 := r2782(19 to 19);
    r2805 := r2782(20 to 20);
    r2806 := r2782(21 to 21);
    r2807 := r2782(22 to 22);
    r2808 := r2782(23 to 23);
    r2809 := r2782(24 to 24);
    r2810 := r2782(25 to 25);
    r2811 := r2782(26 to 26);
    r2812 := r2782(27 to 27);
    r2813 := r2782(28 to 28);
    r2814 := r2782(29 to 29);
    r2815 := r2782(30 to 30);
    r2816 := r2782(31 to 31);
    b2817 := true;
    b2818 := true;
    b2819 := true;
    b2820 := true;
    b2821 := true;
    b2822 := true;
    b2823 := true;
    b2824 := true;
    b2825 := true;
    b2826 := true;
    b2827 := true;
    b2828 := true;
    b2829 := true;
    b2830 := true;
    b2831 := true;
    b2832 := true;
    b2833 := true;
    b2834 := true;
    b2835 := true;
    b2836 := true;
    b2837 := true;
    b2838 := true;
    b2839 := true;
    b2840 := true;
    b2841 := true;
    b2842 := true;
    b2843 := true;
    b2844 := true;
    b2845 := true;
    b2846 := true;
    b2847 := true;
    b2848 := true;
    b2849 := (b2784 AND (b2817 AND (b2818 AND (b2819 AND (b2820 AND (b2821 AND (b2822 AND (b2823 AND (b2824 AND (b2825 AND (b2826 AND (b2827 AND (b2828 AND (b2829 AND (b2830 AND (b2831 AND (b2832 AND (b2833 AND (b2834 AND (b2835 AND (b2836 AND (b2837 AND (b2838 AND (b2839 AND (b2840 AND (b2841 AND (b2842 AND (b2843 AND (b2844 AND (b2845 AND (b2846 AND (b2847 AND b2848))))))))))))))))))))))))))))))));
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    r2850 := (r2795 & r2796 & r2797 & r2798 & r2799 & r2800 & r2801 & r2802 & r2803 & r2804 & r2805 & r2806 & r2807 & r2808 & r2809 & r2810 & r2811 & r2812 & r2813 & r2814 & r2815 & r2816 & r2785 & r2786 & r2787 & r2788 & r2789 & r2790 & r2791 & r2792 & r2793 & r2794);
    r2783 := r2850;
    return r2783;
  end rewire_RWPreluderotateR22_2781;
  function rewire_RWPreluderotateR13_2709(r2710 : std_logic_vector) return std_logic_vector
  is
    variable r2778 : std_logic_vector(0 to 31) := (others => '0');
    variable b2777 : boolean := false;
    variable b2776 : boolean := false;
    variable b2775 : boolean := false;
    variable b2774 : boolean := false;
    variable b2773 : boolean := false;
    variable b2772 : boolean := false;
    variable b2771 : boolean := false;
    variable b2770 : boolean := false;
    variable b2769 : boolean := false;
    variable b2768 : boolean := false;
    variable b2767 : boolean := false;
    variable b2766 : boolean := false;
    variable b2765 : boolean := false;
    variable b2764 : boolean := false;
    variable b2763 : boolean := false;
    variable b2762 : boolean := false;
    variable b2761 : boolean := false;
    variable b2760 : boolean := false;
    variable b2759 : boolean := false;
    variable b2758 : boolean := false;
    variable b2757 : boolean := false;
    variable b2756 : boolean := false;
    variable b2755 : boolean := false;
    variable b2754 : boolean := false;
    variable b2753 : boolean := false;
    variable b2752 : boolean := false;
    variable b2751 : boolean := false;
    variable b2750 : boolean := false;
    variable b2749 : boolean := false;
    variable b2748 : boolean := false;
    variable b2747 : boolean := false;
    variable b2746 : boolean := false;
    variable b2745 : boolean := false;
    variable r2744 : std_logic_vector(0 to 0) := (others => '0');
    variable r2743 : std_logic_vector(0 to 0) := (others => '0');
    variable r2742 : std_logic_vector(0 to 0) := (others => '0');
    variable r2741 : std_logic_vector(0 to 0) := (others => '0');
    variable r2740 : std_logic_vector(0 to 0) := (others => '0');
    variable r2739 : std_logic_vector(0 to 0) := (others => '0');
    variable r2738 : std_logic_vector(0 to 0) := (others => '0');
    variable r2737 : std_logic_vector(0 to 0) := (others => '0');
    variable r2736 : std_logic_vector(0 to 0) := (others => '0');
    variable r2735 : std_logic_vector(0 to 0) := (others => '0');
    variable r2734 : std_logic_vector(0 to 0) := (others => '0');
    variable r2733 : std_logic_vector(0 to 0) := (others => '0');
    variable r2732 : std_logic_vector(0 to 0) := (others => '0');
    variable r2731 : std_logic_vector(0 to 0) := (others => '0');
    variable r2730 : std_logic_vector(0 to 0) := (others => '0');
    variable r2729 : std_logic_vector(0 to 0) := (others => '0');
    variable r2728 : std_logic_vector(0 to 0) := (others => '0');
    variable r2727 : std_logic_vector(0 to 0) := (others => '0');
    variable r2726 : std_logic_vector(0 to 0) := (others => '0');
    variable r2725 : std_logic_vector(0 to 0) := (others => '0');
    variable r2724 : std_logic_vector(0 to 0) := (others => '0');
    variable r2723 : std_logic_vector(0 to 0) := (others => '0');
    variable r2722 : std_logic_vector(0 to 0) := (others => '0');
    variable r2721 : std_logic_vector(0 to 0) := (others => '0');
    variable r2720 : std_logic_vector(0 to 0) := (others => '0');
    variable r2719 : std_logic_vector(0 to 0) := (others => '0');
    variable r2718 : std_logic_vector(0 to 0) := (others => '0');
    variable r2717 : std_logic_vector(0 to 0) := (others => '0');
    variable r2716 : std_logic_vector(0 to 0) := (others => '0');
    variable r2715 : std_logic_vector(0 to 0) := (others => '0');
    variable r2714 : std_logic_vector(0 to 0) := (others => '0');
    variable r2713 : std_logic_vector(0 to 0) := (others => '0');
    variable b2712 : boolean := false;
    variable r2711 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    b2712 := true;
    r2713 := r2710(0 to 0);
    r2714 := r2710(1 to 1);
    r2715 := r2710(2 to 2);
    r2716 := r2710(3 to 3);
    r2717 := r2710(4 to 4);
    r2718 := r2710(5 to 5);
    r2719 := r2710(6 to 6);
    r2720 := r2710(7 to 7);
    r2721 := r2710(8 to 8);
    r2722 := r2710(9 to 9);
    r2723 := r2710(10 to 10);
    r2724 := r2710(11 to 11);
    r2725 := r2710(12 to 12);
    r2726 := r2710(13 to 13);
    r2727 := r2710(14 to 14);
    r2728 := r2710(15 to 15);
    r2729 := r2710(16 to 16);
    r2730 := r2710(17 to 17);
    r2731 := r2710(18 to 18);
    r2732 := r2710(19 to 19);
    r2733 := r2710(20 to 20);
    r2734 := r2710(21 to 21);
    r2735 := r2710(22 to 22);
    r2736 := r2710(23 to 23);
    r2737 := r2710(24 to 24);
    r2738 := r2710(25 to 25);
    r2739 := r2710(26 to 26);
    r2740 := r2710(27 to 27);
    r2741 := r2710(28 to 28);
    r2742 := r2710(29 to 29);
    r2743 := r2710(30 to 30);
    r2744 := r2710(31 to 31);
    b2745 := true;
    b2746 := true;
    b2747 := true;
    b2748 := true;
    b2749 := true;
    b2750 := true;
    b2751 := true;
    b2752 := true;
    b2753 := true;
    b2754 := true;
    b2755 := true;
    b2756 := true;
    b2757 := true;
    b2758 := true;
    b2759 := true;
    b2760 := true;
    b2761 := true;
    b2762 := true;
    b2763 := true;
    b2764 := true;
    b2765 := true;
    b2766 := true;
    b2767 := true;
    b2768 := true;
    b2769 := true;
    b2770 := true;
    b2771 := true;
    b2772 := true;
    b2773 := true;
    b2774 := true;
    b2775 := true;
    b2776 := true;
    b2777 := (b2712 AND (b2745 AND (b2746 AND (b2747 AND (b2748 AND (b2749 AND (b2750 AND (b2751 AND (b2752 AND (b2753 AND (b2754 AND (b2755 AND (b2756 AND (b2757 AND (b2758 AND (b2759 AND (b2760 AND (b2761 AND (b2762 AND (b2763 AND (b2764 AND (b2765 AND (b2766 AND (b2767 AND (b2768 AND (b2769 AND (b2770 AND (b2771 AND (b2772 AND (b2773 AND (b2774 AND (b2775 AND b2776))))))))))))))))))))))))))))))));
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    r2778 := (r2732 & r2733 & r2734 & r2735 & r2736 & r2737 & r2738 & r2739 & r2740 & r2741 & r2742 & r2743 & r2744 & r2713 & r2714 & r2715 & r2716 & r2717 & r2718 & r2719 & r2720 & r2721 & r2722 & r2723 & r2724 & r2725 & r2726 & r2727 & r2728 & r2729 & r2730 & r2731);
    r2711 := r2778;
    return r2711;
  end rewire_RWPreluderotateR13_2709;
  function rewire_RWPreluderotateR2_2638(r2639 : std_logic_vector) return std_logic_vector
  is
    variable r2707 : std_logic_vector(0 to 31) := (others => '0');
    variable b2706 : boolean := false;
    variable b2705 : boolean := false;
    variable b2704 : boolean := false;
    variable b2703 : boolean := false;
    variable b2702 : boolean := false;
    variable b2701 : boolean := false;
    variable b2700 : boolean := false;
    variable b2699 : boolean := false;
    variable b2698 : boolean := false;
    variable b2697 : boolean := false;
    variable b2696 : boolean := false;
    variable b2695 : boolean := false;
    variable b2694 : boolean := false;
    variable b2693 : boolean := false;
    variable b2692 : boolean := false;
    variable b2691 : boolean := false;
    variable b2690 : boolean := false;
    variable b2689 : boolean := false;
    variable b2688 : boolean := false;
    variable b2687 : boolean := false;
    variable b2686 : boolean := false;
    variable b2685 : boolean := false;
    variable b2684 : boolean := false;
    variable b2683 : boolean := false;
    variable b2682 : boolean := false;
    variable b2681 : boolean := false;
    variable b2680 : boolean := false;
    variable b2679 : boolean := false;
    variable b2678 : boolean := false;
    variable b2677 : boolean := false;
    variable b2676 : boolean := false;
    variable b2675 : boolean := false;
    variable b2674 : boolean := false;
    variable r2673 : std_logic_vector(0 to 0) := (others => '0');
    variable r2672 : std_logic_vector(0 to 0) := (others => '0');
    variable r2671 : std_logic_vector(0 to 0) := (others => '0');
    variable r2670 : std_logic_vector(0 to 0) := (others => '0');
    variable r2669 : std_logic_vector(0 to 0) := (others => '0');
    variable r2668 : std_logic_vector(0 to 0) := (others => '0');
    variable r2667 : std_logic_vector(0 to 0) := (others => '0');
    variable r2666 : std_logic_vector(0 to 0) := (others => '0');
    variable r2665 : std_logic_vector(0 to 0) := (others => '0');
    variable r2664 : std_logic_vector(0 to 0) := (others => '0');
    variable r2663 : std_logic_vector(0 to 0) := (others => '0');
    variable r2662 : std_logic_vector(0 to 0) := (others => '0');
    variable r2661 : std_logic_vector(0 to 0) := (others => '0');
    variable r2660 : std_logic_vector(0 to 0) := (others => '0');
    variable r2659 : std_logic_vector(0 to 0) := (others => '0');
    variable r2658 : std_logic_vector(0 to 0) := (others => '0');
    variable r2657 : std_logic_vector(0 to 0) := (others => '0');
    variable r2656 : std_logic_vector(0 to 0) := (others => '0');
    variable r2655 : std_logic_vector(0 to 0) := (others => '0');
    variable r2654 : std_logic_vector(0 to 0) := (others => '0');
    variable r2653 : std_logic_vector(0 to 0) := (others => '0');
    variable r2652 : std_logic_vector(0 to 0) := (others => '0');
    variable r2651 : std_logic_vector(0 to 0) := (others => '0');
    variable r2650 : std_logic_vector(0 to 0) := (others => '0');
    variable r2649 : std_logic_vector(0 to 0) := (others => '0');
    variable r2648 : std_logic_vector(0 to 0) := (others => '0');
    variable r2647 : std_logic_vector(0 to 0) := (others => '0');
    variable r2646 : std_logic_vector(0 to 0) := (others => '0');
    variable r2645 : std_logic_vector(0 to 0) := (others => '0');
    variable r2644 : std_logic_vector(0 to 0) := (others => '0');
    variable r2643 : std_logic_vector(0 to 0) := (others => '0');
    variable r2642 : std_logic_vector(0 to 0) := (others => '0');
    variable b2641 : boolean := false;
    variable r2640 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    b2641 := true;
    r2642 := r2639(0 to 0);
    r2643 := r2639(1 to 1);
    r2644 := r2639(2 to 2);
    r2645 := r2639(3 to 3);
    r2646 := r2639(4 to 4);
    r2647 := r2639(5 to 5);
    r2648 := r2639(6 to 6);
    r2649 := r2639(7 to 7);
    r2650 := r2639(8 to 8);
    r2651 := r2639(9 to 9);
    r2652 := r2639(10 to 10);
    r2653 := r2639(11 to 11);
    r2654 := r2639(12 to 12);
    r2655 := r2639(13 to 13);
    r2656 := r2639(14 to 14);
    r2657 := r2639(15 to 15);
    r2658 := r2639(16 to 16);
    r2659 := r2639(17 to 17);
    r2660 := r2639(18 to 18);
    r2661 := r2639(19 to 19);
    r2662 := r2639(20 to 20);
    r2663 := r2639(21 to 21);
    r2664 := r2639(22 to 22);
    r2665 := r2639(23 to 23);
    r2666 := r2639(24 to 24);
    r2667 := r2639(25 to 25);
    r2668 := r2639(26 to 26);
    r2669 := r2639(27 to 27);
    r2670 := r2639(28 to 28);
    r2671 := r2639(29 to 29);
    r2672 := r2639(30 to 30);
    r2673 := r2639(31 to 31);
    b2674 := true;
    b2675 := true;
    b2676 := true;
    b2677 := true;
    b2678 := true;
    b2679 := true;
    b2680 := true;
    b2681 := true;
    b2682 := true;
    b2683 := true;
    b2684 := true;
    b2685 := true;
    b2686 := true;
    b2687 := true;
    b2688 := true;
    b2689 := true;
    b2690 := true;
    b2691 := true;
    b2692 := true;
    b2693 := true;
    b2694 := true;
    b2695 := true;
    b2696 := true;
    b2697 := true;
    b2698 := true;
    b2699 := true;
    b2700 := true;
    b2701 := true;
    b2702 := true;
    b2703 := true;
    b2704 := true;
    b2705 := true;
    b2706 := (b2641 AND (b2674 AND (b2675 AND (b2676 AND (b2677 AND (b2678 AND (b2679 AND (b2680 AND (b2681 AND (b2682 AND (b2683 AND (b2684 AND (b2685 AND (b2686 AND (b2687 AND (b2688 AND (b2689 AND (b2690 AND (b2691 AND (b2692 AND (b2693 AND (b2694 AND (b2695 AND (b2696 AND (b2697 AND (b2698 AND (b2699 AND (b2700 AND (b2701 AND (b2702 AND (b2703 AND (b2704 AND b2705))))))))))))))))))))))))))))))));
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    r2707 := (r2672 & r2673 & r2642 & r2643 & r2644 & r2645 & r2646 & r2647 & r2648 & r2649 & r2650 & r2651 & r2652 & r2653 & r2654 & r2655 & r2656 & r2657 & r2658 & r2659 & r2660 & r2661 & r2662 & r2663 & r2664 & r2665 & r2666 & r2667 & r2668 & r2669 & r2670 & r2671);
    r2640 := r2707;
    return r2640;
  end rewire_RWPreluderotateR2_2638;
  function rewire_Mainch_2623(r2624 : std_logic_vector ; r2625 : std_logic_vector ; r2626 : std_logic_vector) return std_logic_vector
  is
    variable r2630 : std_logic_vector(0 to 31) := (others => '0');
    variable r2629 : std_logic_vector(0 to 31) := (others => '0');
    variable r2628 : std_logic_vector(0 to 31) := (others => '0');
    variable r2627 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r2627 := w32And(r2624,r2625);
    null;
    r2628 := w32Not(r2624);
    null;
    r2629 := w32And(r2628,r2626);
    r2630 := w32Xor(r2627,r2629);
    return r2630;
  end rewire_Mainch_2623;
  function rewire_Mainbigsigma1_2405(r2406 : std_logic_vector) return std_logic_vector
  is
    variable r2621 : std_logic_vector(0 to 31) := (others => '0');
    variable r2620 : std_logic_vector(0 to 31) := (others => '0');
    variable r2551 : std_logic_vector(0 to 31) := (others => '0');
    variable r2549 : std_logic_vector(0 to 31) := (others => '0');
    variable r2548 : std_logic_vector(0 to 31) := (others => '0');
    variable r2479 : std_logic_vector(0 to 31) := (others => '0');
    variable r2477 : std_logic_vector(0 to 31) := (others => '0');
    variable r2408 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    r2477 := rewire_RWPreluderotateR6_2407(r2406);
    null;
    r2548 := rewire_RWPreluderotateR11_2478(r2406);
    r2549 := w32Xor(r2477,r2548);
    null;
    r2620 := rewire_RWPreluderotateR25_2550(r2406);
    r2621 := w32Xor(r2549,r2620);
    return r2621;
  end rewire_Mainbigsigma1_2405;
  function rewire_RWPreluderotateR25_2550(r2551 : std_logic_vector) return std_logic_vector
  is
    variable r2619 : std_logic_vector(0 to 31) := (others => '0');
    variable b2618 : boolean := false;
    variable b2617 : boolean := false;
    variable b2616 : boolean := false;
    variable b2615 : boolean := false;
    variable b2614 : boolean := false;
    variable b2613 : boolean := false;
    variable b2612 : boolean := false;
    variable b2611 : boolean := false;
    variable b2610 : boolean := false;
    variable b2609 : boolean := false;
    variable b2608 : boolean := false;
    variable b2607 : boolean := false;
    variable b2606 : boolean := false;
    variable b2605 : boolean := false;
    variable b2604 : boolean := false;
    variable b2603 : boolean := false;
    variable b2602 : boolean := false;
    variable b2601 : boolean := false;
    variable b2600 : boolean := false;
    variable b2599 : boolean := false;
    variable b2598 : boolean := false;
    variable b2597 : boolean := false;
    variable b2596 : boolean := false;
    variable b2595 : boolean := false;
    variable b2594 : boolean := false;
    variable b2593 : boolean := false;
    variable b2592 : boolean := false;
    variable b2591 : boolean := false;
    variable b2590 : boolean := false;
    variable b2589 : boolean := false;
    variable b2588 : boolean := false;
    variable b2587 : boolean := false;
    variable b2586 : boolean := false;
    variable r2585 : std_logic_vector(0 to 0) := (others => '0');
    variable r2584 : std_logic_vector(0 to 0) := (others => '0');
    variable r2583 : std_logic_vector(0 to 0) := (others => '0');
    variable r2582 : std_logic_vector(0 to 0) := (others => '0');
    variable r2581 : std_logic_vector(0 to 0) := (others => '0');
    variable r2580 : std_logic_vector(0 to 0) := (others => '0');
    variable r2579 : std_logic_vector(0 to 0) := (others => '0');
    variable r2578 : std_logic_vector(0 to 0) := (others => '0');
    variable r2577 : std_logic_vector(0 to 0) := (others => '0');
    variable r2576 : std_logic_vector(0 to 0) := (others => '0');
    variable r2575 : std_logic_vector(0 to 0) := (others => '0');
    variable r2574 : std_logic_vector(0 to 0) := (others => '0');
    variable r2573 : std_logic_vector(0 to 0) := (others => '0');
    variable r2572 : std_logic_vector(0 to 0) := (others => '0');
    variable r2571 : std_logic_vector(0 to 0) := (others => '0');
    variable r2570 : std_logic_vector(0 to 0) := (others => '0');
    variable r2569 : std_logic_vector(0 to 0) := (others => '0');
    variable r2568 : std_logic_vector(0 to 0) := (others => '0');
    variable r2567 : std_logic_vector(0 to 0) := (others => '0');
    variable r2566 : std_logic_vector(0 to 0) := (others => '0');
    variable r2565 : std_logic_vector(0 to 0) := (others => '0');
    variable r2564 : std_logic_vector(0 to 0) := (others => '0');
    variable r2563 : std_logic_vector(0 to 0) := (others => '0');
    variable r2562 : std_logic_vector(0 to 0) := (others => '0');
    variable r2561 : std_logic_vector(0 to 0) := (others => '0');
    variable r2560 : std_logic_vector(0 to 0) := (others => '0');
    variable r2559 : std_logic_vector(0 to 0) := (others => '0');
    variable r2558 : std_logic_vector(0 to 0) := (others => '0');
    variable r2557 : std_logic_vector(0 to 0) := (others => '0');
    variable r2556 : std_logic_vector(0 to 0) := (others => '0');
    variable r2555 : std_logic_vector(0 to 0) := (others => '0');
    variable r2554 : std_logic_vector(0 to 0) := (others => '0');
    variable b2553 : boolean := false;
    variable r2552 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    b2553 := true;
    r2554 := r2551(0 to 0);
    r2555 := r2551(1 to 1);
    r2556 := r2551(2 to 2);
    r2557 := r2551(3 to 3);
    r2558 := r2551(4 to 4);
    r2559 := r2551(5 to 5);
    r2560 := r2551(6 to 6);
    r2561 := r2551(7 to 7);
    r2562 := r2551(8 to 8);
    r2563 := r2551(9 to 9);
    r2564 := r2551(10 to 10);
    r2565 := r2551(11 to 11);
    r2566 := r2551(12 to 12);
    r2567 := r2551(13 to 13);
    r2568 := r2551(14 to 14);
    r2569 := r2551(15 to 15);
    r2570 := r2551(16 to 16);
    r2571 := r2551(17 to 17);
    r2572 := r2551(18 to 18);
    r2573 := r2551(19 to 19);
    r2574 := r2551(20 to 20);
    r2575 := r2551(21 to 21);
    r2576 := r2551(22 to 22);
    r2577 := r2551(23 to 23);
    r2578 := r2551(24 to 24);
    r2579 := r2551(25 to 25);
    r2580 := r2551(26 to 26);
    r2581 := r2551(27 to 27);
    r2582 := r2551(28 to 28);
    r2583 := r2551(29 to 29);
    r2584 := r2551(30 to 30);
    r2585 := r2551(31 to 31);
    b2586 := true;
    b2587 := true;
    b2588 := true;
    b2589 := true;
    b2590 := true;
    b2591 := true;
    b2592 := true;
    b2593 := true;
    b2594 := true;
    b2595 := true;
    b2596 := true;
    b2597 := true;
    b2598 := true;
    b2599 := true;
    b2600 := true;
    b2601 := true;
    b2602 := true;
    b2603 := true;
    b2604 := true;
    b2605 := true;
    b2606 := true;
    b2607 := true;
    b2608 := true;
    b2609 := true;
    b2610 := true;
    b2611 := true;
    b2612 := true;
    b2613 := true;
    b2614 := true;
    b2615 := true;
    b2616 := true;
    b2617 := true;
    b2618 := (b2553 AND (b2586 AND (b2587 AND (b2588 AND (b2589 AND (b2590 AND (b2591 AND (b2592 AND (b2593 AND (b2594 AND (b2595 AND (b2596 AND (b2597 AND (b2598 AND (b2599 AND (b2600 AND (b2601 AND (b2602 AND (b2603 AND (b2604 AND (b2605 AND (b2606 AND (b2607 AND (b2608 AND (b2609 AND (b2610 AND (b2611 AND (b2612 AND (b2613 AND (b2614 AND (b2615 AND (b2616 AND b2617))))))))))))))))))))))))))))))));
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    r2619 := (r2561 & r2562 & r2563 & r2564 & r2565 & r2566 & r2567 & r2568 & r2569 & r2570 & r2571 & r2572 & r2573 & r2574 & r2575 & r2576 & r2577 & r2578 & r2579 & r2580 & r2581 & r2582 & r2583 & r2584 & r2585 & r2554 & r2555 & r2556 & r2557 & r2558 & r2559 & r2560);
    r2552 := r2619;
    return r2552;
  end rewire_RWPreluderotateR25_2550;
  function rewire_RWPreluderotateR11_2478(r2479 : std_logic_vector) return std_logic_vector
  is
    variable r2547 : std_logic_vector(0 to 31) := (others => '0');
    variable b2546 : boolean := false;
    variable b2545 : boolean := false;
    variable b2544 : boolean := false;
    variable b2543 : boolean := false;
    variable b2542 : boolean := false;
    variable b2541 : boolean := false;
    variable b2540 : boolean := false;
    variable b2539 : boolean := false;
    variable b2538 : boolean := false;
    variable b2537 : boolean := false;
    variable b2536 : boolean := false;
    variable b2535 : boolean := false;
    variable b2534 : boolean := false;
    variable b2533 : boolean := false;
    variable b2532 : boolean := false;
    variable b2531 : boolean := false;
    variable b2530 : boolean := false;
    variable b2529 : boolean := false;
    variable b2528 : boolean := false;
    variable b2527 : boolean := false;
    variable b2526 : boolean := false;
    variable b2525 : boolean := false;
    variable b2524 : boolean := false;
    variable b2523 : boolean := false;
    variable b2522 : boolean := false;
    variable b2521 : boolean := false;
    variable b2520 : boolean := false;
    variable b2519 : boolean := false;
    variable b2518 : boolean := false;
    variable b2517 : boolean := false;
    variable b2516 : boolean := false;
    variable b2515 : boolean := false;
    variable b2514 : boolean := false;
    variable r2513 : std_logic_vector(0 to 0) := (others => '0');
    variable r2512 : std_logic_vector(0 to 0) := (others => '0');
    variable r2511 : std_logic_vector(0 to 0) := (others => '0');
    variable r2510 : std_logic_vector(0 to 0) := (others => '0');
    variable r2509 : std_logic_vector(0 to 0) := (others => '0');
    variable r2508 : std_logic_vector(0 to 0) := (others => '0');
    variable r2507 : std_logic_vector(0 to 0) := (others => '0');
    variable r2506 : std_logic_vector(0 to 0) := (others => '0');
    variable r2505 : std_logic_vector(0 to 0) := (others => '0');
    variable r2504 : std_logic_vector(0 to 0) := (others => '0');
    variable r2503 : std_logic_vector(0 to 0) := (others => '0');
    variable r2502 : std_logic_vector(0 to 0) := (others => '0');
    variable r2501 : std_logic_vector(0 to 0) := (others => '0');
    variable r2500 : std_logic_vector(0 to 0) := (others => '0');
    variable r2499 : std_logic_vector(0 to 0) := (others => '0');
    variable r2498 : std_logic_vector(0 to 0) := (others => '0');
    variable r2497 : std_logic_vector(0 to 0) := (others => '0');
    variable r2496 : std_logic_vector(0 to 0) := (others => '0');
    variable r2495 : std_logic_vector(0 to 0) := (others => '0');
    variable r2494 : std_logic_vector(0 to 0) := (others => '0');
    variable r2493 : std_logic_vector(0 to 0) := (others => '0');
    variable r2492 : std_logic_vector(0 to 0) := (others => '0');
    variable r2491 : std_logic_vector(0 to 0) := (others => '0');
    variable r2490 : std_logic_vector(0 to 0) := (others => '0');
    variable r2489 : std_logic_vector(0 to 0) := (others => '0');
    variable r2488 : std_logic_vector(0 to 0) := (others => '0');
    variable r2487 : std_logic_vector(0 to 0) := (others => '0');
    variable r2486 : std_logic_vector(0 to 0) := (others => '0');
    variable r2485 : std_logic_vector(0 to 0) := (others => '0');
    variable r2484 : std_logic_vector(0 to 0) := (others => '0');
    variable r2483 : std_logic_vector(0 to 0) := (others => '0');
    variable r2482 : std_logic_vector(0 to 0) := (others => '0');
    variable b2481 : boolean := false;
    variable r2480 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    b2481 := true;
    r2482 := r2479(0 to 0);
    r2483 := r2479(1 to 1);
    r2484 := r2479(2 to 2);
    r2485 := r2479(3 to 3);
    r2486 := r2479(4 to 4);
    r2487 := r2479(5 to 5);
    r2488 := r2479(6 to 6);
    r2489 := r2479(7 to 7);
    r2490 := r2479(8 to 8);
    r2491 := r2479(9 to 9);
    r2492 := r2479(10 to 10);
    r2493 := r2479(11 to 11);
    r2494 := r2479(12 to 12);
    r2495 := r2479(13 to 13);
    r2496 := r2479(14 to 14);
    r2497 := r2479(15 to 15);
    r2498 := r2479(16 to 16);
    r2499 := r2479(17 to 17);
    r2500 := r2479(18 to 18);
    r2501 := r2479(19 to 19);
    r2502 := r2479(20 to 20);
    r2503 := r2479(21 to 21);
    r2504 := r2479(22 to 22);
    r2505 := r2479(23 to 23);
    r2506 := r2479(24 to 24);
    r2507 := r2479(25 to 25);
    r2508 := r2479(26 to 26);
    r2509 := r2479(27 to 27);
    r2510 := r2479(28 to 28);
    r2511 := r2479(29 to 29);
    r2512 := r2479(30 to 30);
    r2513 := r2479(31 to 31);
    b2514 := true;
    b2515 := true;
    b2516 := true;
    b2517 := true;
    b2518 := true;
    b2519 := true;
    b2520 := true;
    b2521 := true;
    b2522 := true;
    b2523 := true;
    b2524 := true;
    b2525 := true;
    b2526 := true;
    b2527 := true;
    b2528 := true;
    b2529 := true;
    b2530 := true;
    b2531 := true;
    b2532 := true;
    b2533 := true;
    b2534 := true;
    b2535 := true;
    b2536 := true;
    b2537 := true;
    b2538 := true;
    b2539 := true;
    b2540 := true;
    b2541 := true;
    b2542 := true;
    b2543 := true;
    b2544 := true;
    b2545 := true;
    b2546 := (b2481 AND (b2514 AND (b2515 AND (b2516 AND (b2517 AND (b2518 AND (b2519 AND (b2520 AND (b2521 AND (b2522 AND (b2523 AND (b2524 AND (b2525 AND (b2526 AND (b2527 AND (b2528 AND (b2529 AND (b2530 AND (b2531 AND (b2532 AND (b2533 AND (b2534 AND (b2535 AND (b2536 AND (b2537 AND (b2538 AND (b2539 AND (b2540 AND (b2541 AND (b2542 AND (b2543 AND (b2544 AND b2545))))))))))))))))))))))))))))))));
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    r2547 := (r2503 & r2504 & r2505 & r2506 & r2507 & r2508 & r2509 & r2510 & r2511 & r2512 & r2513 & r2482 & r2483 & r2484 & r2485 & r2486 & r2487 & r2488 & r2489 & r2490 & r2491 & r2492 & r2493 & r2494 & r2495 & r2496 & r2497 & r2498 & r2499 & r2500 & r2501 & r2502);
    r2480 := r2547;
    return r2480;
  end rewire_RWPreluderotateR11_2478;
  function rewire_RWPreluderotateR6_2407(r2408 : std_logic_vector) return std_logic_vector
  is
    variable r2476 : std_logic_vector(0 to 31) := (others => '0');
    variable b2475 : boolean := false;
    variable b2474 : boolean := false;
    variable b2473 : boolean := false;
    variable b2472 : boolean := false;
    variable b2471 : boolean := false;
    variable b2470 : boolean := false;
    variable b2469 : boolean := false;
    variable b2468 : boolean := false;
    variable b2467 : boolean := false;
    variable b2466 : boolean := false;
    variable b2465 : boolean := false;
    variable b2464 : boolean := false;
    variable b2463 : boolean := false;
    variable b2462 : boolean := false;
    variable b2461 : boolean := false;
    variable b2460 : boolean := false;
    variable b2459 : boolean := false;
    variable b2458 : boolean := false;
    variable b2457 : boolean := false;
    variable b2456 : boolean := false;
    variable b2455 : boolean := false;
    variable b2454 : boolean := false;
    variable b2453 : boolean := false;
    variable b2452 : boolean := false;
    variable b2451 : boolean := false;
    variable b2450 : boolean := false;
    variable b2449 : boolean := false;
    variable b2448 : boolean := false;
    variable b2447 : boolean := false;
    variable b2446 : boolean := false;
    variable b2445 : boolean := false;
    variable b2444 : boolean := false;
    variable b2443 : boolean := false;
    variable r2442 : std_logic_vector(0 to 0) := (others => '0');
    variable r2441 : std_logic_vector(0 to 0) := (others => '0');
    variable r2440 : std_logic_vector(0 to 0) := (others => '0');
    variable r2439 : std_logic_vector(0 to 0) := (others => '0');
    variable r2438 : std_logic_vector(0 to 0) := (others => '0');
    variable r2437 : std_logic_vector(0 to 0) := (others => '0');
    variable r2436 : std_logic_vector(0 to 0) := (others => '0');
    variable r2435 : std_logic_vector(0 to 0) := (others => '0');
    variable r2434 : std_logic_vector(0 to 0) := (others => '0');
    variable r2433 : std_logic_vector(0 to 0) := (others => '0');
    variable r2432 : std_logic_vector(0 to 0) := (others => '0');
    variable r2431 : std_logic_vector(0 to 0) := (others => '0');
    variable r2430 : std_logic_vector(0 to 0) := (others => '0');
    variable r2429 : std_logic_vector(0 to 0) := (others => '0');
    variable r2428 : std_logic_vector(0 to 0) := (others => '0');
    variable r2427 : std_logic_vector(0 to 0) := (others => '0');
    variable r2426 : std_logic_vector(0 to 0) := (others => '0');
    variable r2425 : std_logic_vector(0 to 0) := (others => '0');
    variable r2424 : std_logic_vector(0 to 0) := (others => '0');
    variable r2423 : std_logic_vector(0 to 0) := (others => '0');
    variable r2422 : std_logic_vector(0 to 0) := (others => '0');
    variable r2421 : std_logic_vector(0 to 0) := (others => '0');
    variable r2420 : std_logic_vector(0 to 0) := (others => '0');
    variable r2419 : std_logic_vector(0 to 0) := (others => '0');
    variable r2418 : std_logic_vector(0 to 0) := (others => '0');
    variable r2417 : std_logic_vector(0 to 0) := (others => '0');
    variable r2416 : std_logic_vector(0 to 0) := (others => '0');
    variable r2415 : std_logic_vector(0 to 0) := (others => '0');
    variable r2414 : std_logic_vector(0 to 0) := (others => '0');
    variable r2413 : std_logic_vector(0 to 0) := (others => '0');
    variable r2412 : std_logic_vector(0 to 0) := (others => '0');
    variable r2411 : std_logic_vector(0 to 0) := (others => '0');
    variable b2410 : boolean := false;
    variable r2409 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    b2410 := true;
    r2411 := r2408(0 to 0);
    r2412 := r2408(1 to 1);
    r2413 := r2408(2 to 2);
    r2414 := r2408(3 to 3);
    r2415 := r2408(4 to 4);
    r2416 := r2408(5 to 5);
    r2417 := r2408(6 to 6);
    r2418 := r2408(7 to 7);
    r2419 := r2408(8 to 8);
    r2420 := r2408(9 to 9);
    r2421 := r2408(10 to 10);
    r2422 := r2408(11 to 11);
    r2423 := r2408(12 to 12);
    r2424 := r2408(13 to 13);
    r2425 := r2408(14 to 14);
    r2426 := r2408(15 to 15);
    r2427 := r2408(16 to 16);
    r2428 := r2408(17 to 17);
    r2429 := r2408(18 to 18);
    r2430 := r2408(19 to 19);
    r2431 := r2408(20 to 20);
    r2432 := r2408(21 to 21);
    r2433 := r2408(22 to 22);
    r2434 := r2408(23 to 23);
    r2435 := r2408(24 to 24);
    r2436 := r2408(25 to 25);
    r2437 := r2408(26 to 26);
    r2438 := r2408(27 to 27);
    r2439 := r2408(28 to 28);
    r2440 := r2408(29 to 29);
    r2441 := r2408(30 to 30);
    r2442 := r2408(31 to 31);
    b2443 := true;
    b2444 := true;
    b2445 := true;
    b2446 := true;
    b2447 := true;
    b2448 := true;
    b2449 := true;
    b2450 := true;
    b2451 := true;
    b2452 := true;
    b2453 := true;
    b2454 := true;
    b2455 := true;
    b2456 := true;
    b2457 := true;
    b2458 := true;
    b2459 := true;
    b2460 := true;
    b2461 := true;
    b2462 := true;
    b2463 := true;
    b2464 := true;
    b2465 := true;
    b2466 := true;
    b2467 := true;
    b2468 := true;
    b2469 := true;
    b2470 := true;
    b2471 := true;
    b2472 := true;
    b2473 := true;
    b2474 := true;
    b2475 := (b2410 AND (b2443 AND (b2444 AND (b2445 AND (b2446 AND (b2447 AND (b2448 AND (b2449 AND (b2450 AND (b2451 AND (b2452 AND (b2453 AND (b2454 AND (b2455 AND (b2456 AND (b2457 AND (b2458 AND (b2459 AND (b2460 AND (b2461 AND (b2462 AND (b2463 AND (b2464 AND (b2465 AND (b2466 AND (b2467 AND (b2468 AND (b2469 AND (b2470 AND (b2471 AND (b2472 AND (b2473 AND b2474))))))))))))))))))))))))))))))));
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    r2476 := (r2437 & r2438 & r2439 & r2440 & r2441 & r2442 & r2411 & r2412 & r2413 & r2414 & r2415 & r2416 & r2417 & r2418 & r2419 & r2420 & r2421 & r2422 & r2423 & r2424 & r2425 & r2426 & r2427 & r2428 & r2429 & r2430 & r2431 & r2432 & r2433 & r2434 & r2435 & r2436);
    r2409 := r2476;
    return r2409;
  end rewire_RWPreluderotateR6_2407;
  function rewire_MainupdateSched_1861(r1862 : std_logic_vector) return std_logic_vector
  is
    variable r2363 : std_logic_vector(0 to 31) := (others => '0');
    variable r2362 : std_logic_vector(0 to 31) := (others => '0');
    variable r2361 : std_logic_vector(0 to 31) := (others => '0');
    variable r2139 : std_logic_vector(0 to 31) := (others => '0');
    variable r2137 : std_logic_vector(0 to 31) := (others => '0');
    variable r2136 : std_logic_vector(0 to 31) := (others => '0');
    variable r1900 : std_logic_vector(0 to 31) := (others => '0');
    variable r1898 : std_logic_vector(0 to 511) := (others => '0');
    variable b1897 : boolean := false;
    variable b1896 : boolean := false;
    variable b1895 : boolean := false;
    variable b1894 : boolean := false;
    variable b1893 : boolean := false;
    variable b1892 : boolean := false;
    variable b1891 : boolean := false;
    variable b1890 : boolean := false;
    variable b1889 : boolean := false;
    variable b1888 : boolean := false;
    variable b1887 : boolean := false;
    variable b1886 : boolean := false;
    variable b1885 : boolean := false;
    variable b1884 : boolean := false;
    variable b1883 : boolean := false;
    variable b1882 : boolean := false;
    variable b1881 : boolean := false;
    variable r1880 : std_logic_vector(0 to 31) := (others => '0');
    variable r1879 : std_logic_vector(0 to 31) := (others => '0');
    variable r1878 : std_logic_vector(0 to 31) := (others => '0');
    variable r1877 : std_logic_vector(0 to 31) := (others => '0');
    variable r1876 : std_logic_vector(0 to 31) := (others => '0');
    variable r1875 : std_logic_vector(0 to 31) := (others => '0');
    variable r1874 : std_logic_vector(0 to 31) := (others => '0');
    variable r1873 : std_logic_vector(0 to 31) := (others => '0');
    variable r1872 : std_logic_vector(0 to 31) := (others => '0');
    variable r1871 : std_logic_vector(0 to 31) := (others => '0');
    variable r1870 : std_logic_vector(0 to 31) := (others => '0');
    variable r1869 : std_logic_vector(0 to 31) := (others => '0');
    variable r1868 : std_logic_vector(0 to 31) := (others => '0');
    variable r1867 : std_logic_vector(0 to 31) := (others => '0');
    variable r1866 : std_logic_vector(0 to 31) := (others => '0');
    variable r1865 : std_logic_vector(0 to 31) := (others => '0');
    variable b1864 : boolean := false;
    variable r1863 : std_logic_vector(0 to 511) := (others => '0');
  begin
    null;
    b1864 := true;
    r1865 := r1862(0 to 31);
    r1866 := r1862(32 to 63);
    r1867 := r1862(64 to 95);
    r1868 := r1862(96 to 127);
    r1869 := r1862(128 to 159);
    r1870 := r1862(160 to 191);
    r1871 := r1862(192 to 223);
    r1872 := r1862(224 to 255);
    r1873 := r1862(256 to 287);
    r1874 := r1862(288 to 319);
    r1875 := r1862(320 to 351);
    r1876 := r1862(352 to 383);
    r1877 := r1862(384 to 415);
    r1878 := r1862(416 to 447);
    r1879 := r1862(448 to 479);
    r1880 := r1862(480 to 511);
    b1881 := true;
    b1882 := true;
    b1883 := true;
    b1884 := true;
    b1885 := true;
    b1886 := true;
    b1887 := true;
    b1888 := true;
    b1889 := true;
    b1890 := true;
    b1891 := true;
    b1892 := true;
    b1893 := true;
    b1894 := true;
    b1895 := true;
    b1896 := true;
    b1897 := (b1864 AND (b1881 AND (b1882 AND (b1883 AND (b1884 AND (b1885 AND (b1886 AND (b1887 AND (b1888 AND (b1889 AND (b1890 AND (b1891 AND (b1892 AND (b1893 AND (b1894 AND (b1895 AND b1896))))))))))))))));
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    r2136 := rewire_Mainsigma1_1899(r1879);
    null;
    r2137 := w32Plus(r2136,r1874);
    null;
    r2361 := rewire_Mainsigma0_2138(r1866);
    null;
    r2362 := w32Plus(r2361,r1865);
    r2363 := w32Plus(r2137,r2362);
    r1898 := (r1866 & r1867 & r1868 & r1869 & r1870 & r1871 & r1872 & r1873 & r1874 & r1875 & r1876 & r1877 & r1878 & r1879 & r1880 & r2363);
    r1863 := r1898;
    return r1863;
  end rewire_MainupdateSched_1861;
  function rewire_Mainsigma0_2138(r2139 : std_logic_vector) return std_logic_vector
  is
    variable r2360 : std_logic_vector(0 to 31) := (others => '0');
    variable r2359 : std_logic_vector(0 to 31) := (others => '0');
    variable r2284 : std_logic_vector(0 to 31) := (others => '0');
    variable r2282 : std_logic_vector(0 to 31) := (others => '0');
    variable r2281 : std_logic_vector(0 to 31) := (others => '0');
    variable r2212 : std_logic_vector(0 to 31) := (others => '0');
    variable r2210 : std_logic_vector(0 to 31) := (others => '0');
    variable r2141 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    r2210 := rewire_RWPreluderotateR7_2140(r2139);
    null;
    r2281 := rewire_RWPreluderotateR18_2211(r2139);
    r2282 := w32Xor(r2210,r2281);
    null;
    r2359 := rewire_RWPreludeshiftR3_2283(r2139);
    r2360 := w32Xor(r2282,r2359);
    return r2360;
  end rewire_Mainsigma0_2138;
  function rewire_RWPreludeshiftR3_2283(r2284 : std_logic_vector) return std_logic_vector
  is
    variable r2358 : std_logic_vector(0 to 0) := (others => '0');
    variable r2357 : std_logic_vector(0 to 0) := (others => '0');
    variable r2356 : std_logic_vector(0 to 0) := (others => '0');
    variable r2355 : std_logic_vector(0 to 0) := (others => '0');
    variable r2354 : std_logic_vector(0 to 0) := (others => '0');
    variable r2353 : std_logic_vector(0 to 0) := (others => '0');
    variable r2352 : std_logic_vector(0 to 31) := (others => '0');
    variable b2351 : boolean := false;
    variable b2350 : boolean := false;
    variable b2349 : boolean := false;
    variable b2348 : boolean := false;
    variable b2347 : boolean := false;
    variable b2346 : boolean := false;
    variable b2345 : boolean := false;
    variable b2344 : boolean := false;
    variable b2343 : boolean := false;
    variable b2342 : boolean := false;
    variable b2341 : boolean := false;
    variable b2340 : boolean := false;
    variable b2339 : boolean := false;
    variable b2338 : boolean := false;
    variable b2337 : boolean := false;
    variable b2336 : boolean := false;
    variable b2335 : boolean := false;
    variable b2334 : boolean := false;
    variable b2333 : boolean := false;
    variable b2332 : boolean := false;
    variable b2331 : boolean := false;
    variable b2330 : boolean := false;
    variable b2329 : boolean := false;
    variable b2328 : boolean := false;
    variable b2327 : boolean := false;
    variable b2326 : boolean := false;
    variable b2325 : boolean := false;
    variable b2324 : boolean := false;
    variable b2323 : boolean := false;
    variable b2322 : boolean := false;
    variable b2321 : boolean := false;
    variable b2320 : boolean := false;
    variable b2319 : boolean := false;
    variable r2318 : std_logic_vector(0 to 0) := (others => '0');
    variable r2317 : std_logic_vector(0 to 0) := (others => '0');
    variable r2316 : std_logic_vector(0 to 0) := (others => '0');
    variable r2315 : std_logic_vector(0 to 0) := (others => '0');
    variable r2314 : std_logic_vector(0 to 0) := (others => '0');
    variable r2313 : std_logic_vector(0 to 0) := (others => '0');
    variable r2312 : std_logic_vector(0 to 0) := (others => '0');
    variable r2311 : std_logic_vector(0 to 0) := (others => '0');
    variable r2310 : std_logic_vector(0 to 0) := (others => '0');
    variable r2309 : std_logic_vector(0 to 0) := (others => '0');
    variable r2308 : std_logic_vector(0 to 0) := (others => '0');
    variable r2307 : std_logic_vector(0 to 0) := (others => '0');
    variable r2306 : std_logic_vector(0 to 0) := (others => '0');
    variable r2305 : std_logic_vector(0 to 0) := (others => '0');
    variable r2304 : std_logic_vector(0 to 0) := (others => '0');
    variable r2303 : std_logic_vector(0 to 0) := (others => '0');
    variable r2302 : std_logic_vector(0 to 0) := (others => '0');
    variable r2301 : std_logic_vector(0 to 0) := (others => '0');
    variable r2300 : std_logic_vector(0 to 0) := (others => '0');
    variable r2299 : std_logic_vector(0 to 0) := (others => '0');
    variable r2298 : std_logic_vector(0 to 0) := (others => '0');
    variable r2297 : std_logic_vector(0 to 0) := (others => '0');
    variable r2296 : std_logic_vector(0 to 0) := (others => '0');
    variable r2295 : std_logic_vector(0 to 0) := (others => '0');
    variable r2294 : std_logic_vector(0 to 0) := (others => '0');
    variable r2293 : std_logic_vector(0 to 0) := (others => '0');
    variable r2292 : std_logic_vector(0 to 0) := (others => '0');
    variable r2291 : std_logic_vector(0 to 0) := (others => '0');
    variable r2290 : std_logic_vector(0 to 0) := (others => '0');
    variable r2289 : std_logic_vector(0 to 0) := (others => '0');
    variable r2288 : std_logic_vector(0 to 0) := (others => '0');
    variable r2287 : std_logic_vector(0 to 0) := (others => '0');
    variable b2286 : boolean := false;
    variable r2285 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    b2286 := true;
    r2287 := r2284(0 to 0);
    r2288 := r2284(1 to 1);
    r2289 := r2284(2 to 2);
    r2290 := r2284(3 to 3);
    r2291 := r2284(4 to 4);
    r2292 := r2284(5 to 5);
    r2293 := r2284(6 to 6);
    r2294 := r2284(7 to 7);
    r2295 := r2284(8 to 8);
    r2296 := r2284(9 to 9);
    r2297 := r2284(10 to 10);
    r2298 := r2284(11 to 11);
    r2299 := r2284(12 to 12);
    r2300 := r2284(13 to 13);
    r2301 := r2284(14 to 14);
    r2302 := r2284(15 to 15);
    r2303 := r2284(16 to 16);
    r2304 := r2284(17 to 17);
    r2305 := r2284(18 to 18);
    r2306 := r2284(19 to 19);
    r2307 := r2284(20 to 20);
    r2308 := r2284(21 to 21);
    r2309 := r2284(22 to 22);
    r2310 := r2284(23 to 23);
    r2311 := r2284(24 to 24);
    r2312 := r2284(25 to 25);
    r2313 := r2284(26 to 26);
    r2314 := r2284(27 to 27);
    r2315 := r2284(28 to 28);
    r2316 := r2284(29 to 29);
    r2317 := r2284(30 to 30);
    r2318 := r2284(31 to 31);
    b2319 := true;
    b2320 := true;
    b2321 := true;
    b2322 := true;
    b2323 := true;
    b2324 := true;
    b2325 := true;
    b2326 := true;
    b2327 := true;
    b2328 := true;
    b2329 := true;
    b2330 := true;
    b2331 := true;
    b2332 := true;
    b2333 := true;
    b2334 := true;
    b2335 := true;
    b2336 := true;
    b2337 := true;
    b2338 := true;
    b2339 := true;
    b2340 := true;
    b2341 := true;
    b2342 := true;
    b2343 := true;
    b2344 := true;
    b2345 := true;
    b2346 := true;
    b2347 := true;
    b2348 := true;
    b2349 := true;
    b2350 := true;
    b2351 := (b2286 AND (b2319 AND (b2320 AND (b2321 AND (b2322 AND (b2323 AND (b2324 AND (b2325 AND (b2326 AND (b2327 AND (b2328 AND (b2329 AND (b2330 AND (b2331 AND (b2332 AND (b2333 AND (b2334 AND (b2335 AND (b2336 AND (b2337 AND (b2338 AND (b2339 AND (b2340 AND (b2341 AND (b2342 AND (b2343 AND (b2344 AND (b2345 AND (b2346 AND (b2347 AND (b2348 AND (b2349 AND b2350))))))))))))))))))))))))))))))));
    null;
    null;
    r2353 := "0";
    null;
    r2354 := (r2353);
    r2355 := "0";
    null;
    r2356 := (r2355);
    r2357 := "0";
    null;
    r2358 := (r2357);
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    r2352 := (r2354 & r2356 & r2358 & r2287 & r2288 & r2289 & r2290 & r2291 & r2292 & r2293 & r2294 & r2295 & r2296 & r2297 & r2298 & r2299 & r2300 & r2301 & r2302 & r2303 & r2304 & r2305 & r2306 & r2307 & r2308 & r2309 & r2310 & r2311 & r2312 & r2313 & r2314 & r2315);
    r2285 := r2352;
    return r2285;
  end rewire_RWPreludeshiftR3_2283;
  function rewire_RWPreluderotateR18_2211(r2212 : std_logic_vector) return std_logic_vector
  is
    variable r2280 : std_logic_vector(0 to 31) := (others => '0');
    variable b2279 : boolean := false;
    variable b2278 : boolean := false;
    variable b2277 : boolean := false;
    variable b2276 : boolean := false;
    variable b2275 : boolean := false;
    variable b2274 : boolean := false;
    variable b2273 : boolean := false;
    variable b2272 : boolean := false;
    variable b2271 : boolean := false;
    variable b2270 : boolean := false;
    variable b2269 : boolean := false;
    variable b2268 : boolean := false;
    variable b2267 : boolean := false;
    variable b2266 : boolean := false;
    variable b2265 : boolean := false;
    variable b2264 : boolean := false;
    variable b2263 : boolean := false;
    variable b2262 : boolean := false;
    variable b2261 : boolean := false;
    variable b2260 : boolean := false;
    variable b2259 : boolean := false;
    variable b2258 : boolean := false;
    variable b2257 : boolean := false;
    variable b2256 : boolean := false;
    variable b2255 : boolean := false;
    variable b2254 : boolean := false;
    variable b2253 : boolean := false;
    variable b2252 : boolean := false;
    variable b2251 : boolean := false;
    variable b2250 : boolean := false;
    variable b2249 : boolean := false;
    variable b2248 : boolean := false;
    variable b2247 : boolean := false;
    variable r2246 : std_logic_vector(0 to 0) := (others => '0');
    variable r2245 : std_logic_vector(0 to 0) := (others => '0');
    variable r2244 : std_logic_vector(0 to 0) := (others => '0');
    variable r2243 : std_logic_vector(0 to 0) := (others => '0');
    variable r2242 : std_logic_vector(0 to 0) := (others => '0');
    variable r2241 : std_logic_vector(0 to 0) := (others => '0');
    variable r2240 : std_logic_vector(0 to 0) := (others => '0');
    variable r2239 : std_logic_vector(0 to 0) := (others => '0');
    variable r2238 : std_logic_vector(0 to 0) := (others => '0');
    variable r2237 : std_logic_vector(0 to 0) := (others => '0');
    variable r2236 : std_logic_vector(0 to 0) := (others => '0');
    variable r2235 : std_logic_vector(0 to 0) := (others => '0');
    variable r2234 : std_logic_vector(0 to 0) := (others => '0');
    variable r2233 : std_logic_vector(0 to 0) := (others => '0');
    variable r2232 : std_logic_vector(0 to 0) := (others => '0');
    variable r2231 : std_logic_vector(0 to 0) := (others => '0');
    variable r2230 : std_logic_vector(0 to 0) := (others => '0');
    variable r2229 : std_logic_vector(0 to 0) := (others => '0');
    variable r2228 : std_logic_vector(0 to 0) := (others => '0');
    variable r2227 : std_logic_vector(0 to 0) := (others => '0');
    variable r2226 : std_logic_vector(0 to 0) := (others => '0');
    variable r2225 : std_logic_vector(0 to 0) := (others => '0');
    variable r2224 : std_logic_vector(0 to 0) := (others => '0');
    variable r2223 : std_logic_vector(0 to 0) := (others => '0');
    variable r2222 : std_logic_vector(0 to 0) := (others => '0');
    variable r2221 : std_logic_vector(0 to 0) := (others => '0');
    variable r2220 : std_logic_vector(0 to 0) := (others => '0');
    variable r2219 : std_logic_vector(0 to 0) := (others => '0');
    variable r2218 : std_logic_vector(0 to 0) := (others => '0');
    variable r2217 : std_logic_vector(0 to 0) := (others => '0');
    variable r2216 : std_logic_vector(0 to 0) := (others => '0');
    variable r2215 : std_logic_vector(0 to 0) := (others => '0');
    variable b2214 : boolean := false;
    variable r2213 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    b2214 := true;
    r2215 := r2212(0 to 0);
    r2216 := r2212(1 to 1);
    r2217 := r2212(2 to 2);
    r2218 := r2212(3 to 3);
    r2219 := r2212(4 to 4);
    r2220 := r2212(5 to 5);
    r2221 := r2212(6 to 6);
    r2222 := r2212(7 to 7);
    r2223 := r2212(8 to 8);
    r2224 := r2212(9 to 9);
    r2225 := r2212(10 to 10);
    r2226 := r2212(11 to 11);
    r2227 := r2212(12 to 12);
    r2228 := r2212(13 to 13);
    r2229 := r2212(14 to 14);
    r2230 := r2212(15 to 15);
    r2231 := r2212(16 to 16);
    r2232 := r2212(17 to 17);
    r2233 := r2212(18 to 18);
    r2234 := r2212(19 to 19);
    r2235 := r2212(20 to 20);
    r2236 := r2212(21 to 21);
    r2237 := r2212(22 to 22);
    r2238 := r2212(23 to 23);
    r2239 := r2212(24 to 24);
    r2240 := r2212(25 to 25);
    r2241 := r2212(26 to 26);
    r2242 := r2212(27 to 27);
    r2243 := r2212(28 to 28);
    r2244 := r2212(29 to 29);
    r2245 := r2212(30 to 30);
    r2246 := r2212(31 to 31);
    b2247 := true;
    b2248 := true;
    b2249 := true;
    b2250 := true;
    b2251 := true;
    b2252 := true;
    b2253 := true;
    b2254 := true;
    b2255 := true;
    b2256 := true;
    b2257 := true;
    b2258 := true;
    b2259 := true;
    b2260 := true;
    b2261 := true;
    b2262 := true;
    b2263 := true;
    b2264 := true;
    b2265 := true;
    b2266 := true;
    b2267 := true;
    b2268 := true;
    b2269 := true;
    b2270 := true;
    b2271 := true;
    b2272 := true;
    b2273 := true;
    b2274 := true;
    b2275 := true;
    b2276 := true;
    b2277 := true;
    b2278 := true;
    b2279 := (b2214 AND (b2247 AND (b2248 AND (b2249 AND (b2250 AND (b2251 AND (b2252 AND (b2253 AND (b2254 AND (b2255 AND (b2256 AND (b2257 AND (b2258 AND (b2259 AND (b2260 AND (b2261 AND (b2262 AND (b2263 AND (b2264 AND (b2265 AND (b2266 AND (b2267 AND (b2268 AND (b2269 AND (b2270 AND (b2271 AND (b2272 AND (b2273 AND (b2274 AND (b2275 AND (b2276 AND (b2277 AND b2278))))))))))))))))))))))))))))))));
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    r2280 := (r2229 & r2230 & r2231 & r2232 & r2233 & r2234 & r2235 & r2236 & r2237 & r2238 & r2239 & r2240 & r2241 & r2242 & r2243 & r2244 & r2245 & r2246 & r2215 & r2216 & r2217 & r2218 & r2219 & r2220 & r2221 & r2222 & r2223 & r2224 & r2225 & r2226 & r2227 & r2228);
    r2213 := r2280;
    return r2213;
  end rewire_RWPreluderotateR18_2211;
  function rewire_RWPreluderotateR7_2140(r2141 : std_logic_vector) return std_logic_vector
  is
    variable r2209 : std_logic_vector(0 to 31) := (others => '0');
    variable b2208 : boolean := false;
    variable b2207 : boolean := false;
    variable b2206 : boolean := false;
    variable b2205 : boolean := false;
    variable b2204 : boolean := false;
    variable b2203 : boolean := false;
    variable b2202 : boolean := false;
    variable b2201 : boolean := false;
    variable b2200 : boolean := false;
    variable b2199 : boolean := false;
    variable b2198 : boolean := false;
    variable b2197 : boolean := false;
    variable b2196 : boolean := false;
    variable b2195 : boolean := false;
    variable b2194 : boolean := false;
    variable b2193 : boolean := false;
    variable b2192 : boolean := false;
    variable b2191 : boolean := false;
    variable b2190 : boolean := false;
    variable b2189 : boolean := false;
    variable b2188 : boolean := false;
    variable b2187 : boolean := false;
    variable b2186 : boolean := false;
    variable b2185 : boolean := false;
    variable b2184 : boolean := false;
    variable b2183 : boolean := false;
    variable b2182 : boolean := false;
    variable b2181 : boolean := false;
    variable b2180 : boolean := false;
    variable b2179 : boolean := false;
    variable b2178 : boolean := false;
    variable b2177 : boolean := false;
    variable b2176 : boolean := false;
    variable r2175 : std_logic_vector(0 to 0) := (others => '0');
    variable r2174 : std_logic_vector(0 to 0) := (others => '0');
    variable r2173 : std_logic_vector(0 to 0) := (others => '0');
    variable r2172 : std_logic_vector(0 to 0) := (others => '0');
    variable r2171 : std_logic_vector(0 to 0) := (others => '0');
    variable r2170 : std_logic_vector(0 to 0) := (others => '0');
    variable r2169 : std_logic_vector(0 to 0) := (others => '0');
    variable r2168 : std_logic_vector(0 to 0) := (others => '0');
    variable r2167 : std_logic_vector(0 to 0) := (others => '0');
    variable r2166 : std_logic_vector(0 to 0) := (others => '0');
    variable r2165 : std_logic_vector(0 to 0) := (others => '0');
    variable r2164 : std_logic_vector(0 to 0) := (others => '0');
    variable r2163 : std_logic_vector(0 to 0) := (others => '0');
    variable r2162 : std_logic_vector(0 to 0) := (others => '0');
    variable r2161 : std_logic_vector(0 to 0) := (others => '0');
    variable r2160 : std_logic_vector(0 to 0) := (others => '0');
    variable r2159 : std_logic_vector(0 to 0) := (others => '0');
    variable r2158 : std_logic_vector(0 to 0) := (others => '0');
    variable r2157 : std_logic_vector(0 to 0) := (others => '0');
    variable r2156 : std_logic_vector(0 to 0) := (others => '0');
    variable r2155 : std_logic_vector(0 to 0) := (others => '0');
    variable r2154 : std_logic_vector(0 to 0) := (others => '0');
    variable r2153 : std_logic_vector(0 to 0) := (others => '0');
    variable r2152 : std_logic_vector(0 to 0) := (others => '0');
    variable r2151 : std_logic_vector(0 to 0) := (others => '0');
    variable r2150 : std_logic_vector(0 to 0) := (others => '0');
    variable r2149 : std_logic_vector(0 to 0) := (others => '0');
    variable r2148 : std_logic_vector(0 to 0) := (others => '0');
    variable r2147 : std_logic_vector(0 to 0) := (others => '0');
    variable r2146 : std_logic_vector(0 to 0) := (others => '0');
    variable r2145 : std_logic_vector(0 to 0) := (others => '0');
    variable r2144 : std_logic_vector(0 to 0) := (others => '0');
    variable b2143 : boolean := false;
    variable r2142 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    b2143 := true;
    r2144 := r2141(0 to 0);
    r2145 := r2141(1 to 1);
    r2146 := r2141(2 to 2);
    r2147 := r2141(3 to 3);
    r2148 := r2141(4 to 4);
    r2149 := r2141(5 to 5);
    r2150 := r2141(6 to 6);
    r2151 := r2141(7 to 7);
    r2152 := r2141(8 to 8);
    r2153 := r2141(9 to 9);
    r2154 := r2141(10 to 10);
    r2155 := r2141(11 to 11);
    r2156 := r2141(12 to 12);
    r2157 := r2141(13 to 13);
    r2158 := r2141(14 to 14);
    r2159 := r2141(15 to 15);
    r2160 := r2141(16 to 16);
    r2161 := r2141(17 to 17);
    r2162 := r2141(18 to 18);
    r2163 := r2141(19 to 19);
    r2164 := r2141(20 to 20);
    r2165 := r2141(21 to 21);
    r2166 := r2141(22 to 22);
    r2167 := r2141(23 to 23);
    r2168 := r2141(24 to 24);
    r2169 := r2141(25 to 25);
    r2170 := r2141(26 to 26);
    r2171 := r2141(27 to 27);
    r2172 := r2141(28 to 28);
    r2173 := r2141(29 to 29);
    r2174 := r2141(30 to 30);
    r2175 := r2141(31 to 31);
    b2176 := true;
    b2177 := true;
    b2178 := true;
    b2179 := true;
    b2180 := true;
    b2181 := true;
    b2182 := true;
    b2183 := true;
    b2184 := true;
    b2185 := true;
    b2186 := true;
    b2187 := true;
    b2188 := true;
    b2189 := true;
    b2190 := true;
    b2191 := true;
    b2192 := true;
    b2193 := true;
    b2194 := true;
    b2195 := true;
    b2196 := true;
    b2197 := true;
    b2198 := true;
    b2199 := true;
    b2200 := true;
    b2201 := true;
    b2202 := true;
    b2203 := true;
    b2204 := true;
    b2205 := true;
    b2206 := true;
    b2207 := true;
    b2208 := (b2143 AND (b2176 AND (b2177 AND (b2178 AND (b2179 AND (b2180 AND (b2181 AND (b2182 AND (b2183 AND (b2184 AND (b2185 AND (b2186 AND (b2187 AND (b2188 AND (b2189 AND (b2190 AND (b2191 AND (b2192 AND (b2193 AND (b2194 AND (b2195 AND (b2196 AND (b2197 AND (b2198 AND (b2199 AND (b2200 AND (b2201 AND (b2202 AND (b2203 AND (b2204 AND (b2205 AND (b2206 AND b2207))))))))))))))))))))))))))))))));
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    r2209 := (r2169 & r2170 & r2171 & r2172 & r2173 & r2174 & r2175 & r2144 & r2145 & r2146 & r2147 & r2148 & r2149 & r2150 & r2151 & r2152 & r2153 & r2154 & r2155 & r2156 & r2157 & r2158 & r2159 & r2160 & r2161 & r2162 & r2163 & r2164 & r2165 & r2166 & r2167 & r2168);
    r2142 := r2209;
    return r2142;
  end rewire_RWPreluderotateR7_2140;
  function rewire_Mainsigma1_1899(r1900 : std_logic_vector) return std_logic_vector
  is
    variable r2135 : std_logic_vector(0 to 31) := (others => '0');
    variable r2134 : std_logic_vector(0 to 31) := (others => '0');
    variable r2045 : std_logic_vector(0 to 31) := (others => '0');
    variable r2043 : std_logic_vector(0 to 31) := (others => '0');
    variable r2042 : std_logic_vector(0 to 31) := (others => '0');
    variable r1973 : std_logic_vector(0 to 31) := (others => '0');
    variable r1971 : std_logic_vector(0 to 31) := (others => '0');
    variable r1902 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    r1971 := rewire_RWPreluderotateR17_1901(r1900);
    null;
    r2042 := rewire_RWPreluderotateR19_1972(r1900);
    r2043 := w32Xor(r1971,r2042);
    null;
    r2134 := rewire_RWPreludeshiftR10_2044(r1900);
    r2135 := w32Xor(r2043,r2134);
    return r2135;
  end rewire_Mainsigma1_1899;
  function rewire_RWPreludeshiftR10_2044(r2045 : std_logic_vector) return std_logic_vector
  is
    variable r2133 : std_logic_vector(0 to 0) := (others => '0');
    variable r2132 : std_logic_vector(0 to 0) := (others => '0');
    variable r2131 : std_logic_vector(0 to 0) := (others => '0');
    variable r2130 : std_logic_vector(0 to 0) := (others => '0');
    variable r2129 : std_logic_vector(0 to 0) := (others => '0');
    variable r2128 : std_logic_vector(0 to 0) := (others => '0');
    variable r2127 : std_logic_vector(0 to 0) := (others => '0');
    variable r2126 : std_logic_vector(0 to 0) := (others => '0');
    variable r2125 : std_logic_vector(0 to 0) := (others => '0');
    variable r2124 : std_logic_vector(0 to 0) := (others => '0');
    variable r2123 : std_logic_vector(0 to 0) := (others => '0');
    variable r2122 : std_logic_vector(0 to 0) := (others => '0');
    variable r2121 : std_logic_vector(0 to 0) := (others => '0');
    variable r2120 : std_logic_vector(0 to 0) := (others => '0');
    variable r2119 : std_logic_vector(0 to 0) := (others => '0');
    variable r2118 : std_logic_vector(0 to 0) := (others => '0');
    variable r2117 : std_logic_vector(0 to 0) := (others => '0');
    variable r2116 : std_logic_vector(0 to 0) := (others => '0');
    variable r2115 : std_logic_vector(0 to 0) := (others => '0');
    variable r2114 : std_logic_vector(0 to 0) := (others => '0');
    variable r2113 : std_logic_vector(0 to 31) := (others => '0');
    variable b2112 : boolean := false;
    variable b2111 : boolean := false;
    variable b2110 : boolean := false;
    variable b2109 : boolean := false;
    variable b2108 : boolean := false;
    variable b2107 : boolean := false;
    variable b2106 : boolean := false;
    variable b2105 : boolean := false;
    variable b2104 : boolean := false;
    variable b2103 : boolean := false;
    variable b2102 : boolean := false;
    variable b2101 : boolean := false;
    variable b2100 : boolean := false;
    variable b2099 : boolean := false;
    variable b2098 : boolean := false;
    variable b2097 : boolean := false;
    variable b2096 : boolean := false;
    variable b2095 : boolean := false;
    variable b2094 : boolean := false;
    variable b2093 : boolean := false;
    variable b2092 : boolean := false;
    variable b2091 : boolean := false;
    variable b2090 : boolean := false;
    variable b2089 : boolean := false;
    variable b2088 : boolean := false;
    variable b2087 : boolean := false;
    variable b2086 : boolean := false;
    variable b2085 : boolean := false;
    variable b2084 : boolean := false;
    variable b2083 : boolean := false;
    variable b2082 : boolean := false;
    variable b2081 : boolean := false;
    variable b2080 : boolean := false;
    variable r2079 : std_logic_vector(0 to 0) := (others => '0');
    variable r2078 : std_logic_vector(0 to 0) := (others => '0');
    variable r2077 : std_logic_vector(0 to 0) := (others => '0');
    variable r2076 : std_logic_vector(0 to 0) := (others => '0');
    variable r2075 : std_logic_vector(0 to 0) := (others => '0');
    variable r2074 : std_logic_vector(0 to 0) := (others => '0');
    variable r2073 : std_logic_vector(0 to 0) := (others => '0');
    variable r2072 : std_logic_vector(0 to 0) := (others => '0');
    variable r2071 : std_logic_vector(0 to 0) := (others => '0');
    variable r2070 : std_logic_vector(0 to 0) := (others => '0');
    variable r2069 : std_logic_vector(0 to 0) := (others => '0');
    variable r2068 : std_logic_vector(0 to 0) := (others => '0');
    variable r2067 : std_logic_vector(0 to 0) := (others => '0');
    variable r2066 : std_logic_vector(0 to 0) := (others => '0');
    variable r2065 : std_logic_vector(0 to 0) := (others => '0');
    variable r2064 : std_logic_vector(0 to 0) := (others => '0');
    variable r2063 : std_logic_vector(0 to 0) := (others => '0');
    variable r2062 : std_logic_vector(0 to 0) := (others => '0');
    variable r2061 : std_logic_vector(0 to 0) := (others => '0');
    variable r2060 : std_logic_vector(0 to 0) := (others => '0');
    variable r2059 : std_logic_vector(0 to 0) := (others => '0');
    variable r2058 : std_logic_vector(0 to 0) := (others => '0');
    variable r2057 : std_logic_vector(0 to 0) := (others => '0');
    variable r2056 : std_logic_vector(0 to 0) := (others => '0');
    variable r2055 : std_logic_vector(0 to 0) := (others => '0');
    variable r2054 : std_logic_vector(0 to 0) := (others => '0');
    variable r2053 : std_logic_vector(0 to 0) := (others => '0');
    variable r2052 : std_logic_vector(0 to 0) := (others => '0');
    variable r2051 : std_logic_vector(0 to 0) := (others => '0');
    variable r2050 : std_logic_vector(0 to 0) := (others => '0');
    variable r2049 : std_logic_vector(0 to 0) := (others => '0');
    variable r2048 : std_logic_vector(0 to 0) := (others => '0');
    variable b2047 : boolean := false;
    variable r2046 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    b2047 := true;
    r2048 := r2045(0 to 0);
    r2049 := r2045(1 to 1);
    r2050 := r2045(2 to 2);
    r2051 := r2045(3 to 3);
    r2052 := r2045(4 to 4);
    r2053 := r2045(5 to 5);
    r2054 := r2045(6 to 6);
    r2055 := r2045(7 to 7);
    r2056 := r2045(8 to 8);
    r2057 := r2045(9 to 9);
    r2058 := r2045(10 to 10);
    r2059 := r2045(11 to 11);
    r2060 := r2045(12 to 12);
    r2061 := r2045(13 to 13);
    r2062 := r2045(14 to 14);
    r2063 := r2045(15 to 15);
    r2064 := r2045(16 to 16);
    r2065 := r2045(17 to 17);
    r2066 := r2045(18 to 18);
    r2067 := r2045(19 to 19);
    r2068 := r2045(20 to 20);
    r2069 := r2045(21 to 21);
    r2070 := r2045(22 to 22);
    r2071 := r2045(23 to 23);
    r2072 := r2045(24 to 24);
    r2073 := r2045(25 to 25);
    r2074 := r2045(26 to 26);
    r2075 := r2045(27 to 27);
    r2076 := r2045(28 to 28);
    r2077 := r2045(29 to 29);
    r2078 := r2045(30 to 30);
    r2079 := r2045(31 to 31);
    b2080 := true;
    b2081 := true;
    b2082 := true;
    b2083 := true;
    b2084 := true;
    b2085 := true;
    b2086 := true;
    b2087 := true;
    b2088 := true;
    b2089 := true;
    b2090 := true;
    b2091 := true;
    b2092 := true;
    b2093 := true;
    b2094 := true;
    b2095 := true;
    b2096 := true;
    b2097 := true;
    b2098 := true;
    b2099 := true;
    b2100 := true;
    b2101 := true;
    b2102 := true;
    b2103 := true;
    b2104 := true;
    b2105 := true;
    b2106 := true;
    b2107 := true;
    b2108 := true;
    b2109 := true;
    b2110 := true;
    b2111 := true;
    b2112 := (b2047 AND (b2080 AND (b2081 AND (b2082 AND (b2083 AND (b2084 AND (b2085 AND (b2086 AND (b2087 AND (b2088 AND (b2089 AND (b2090 AND (b2091 AND (b2092 AND (b2093 AND (b2094 AND (b2095 AND (b2096 AND (b2097 AND (b2098 AND (b2099 AND (b2100 AND (b2101 AND (b2102 AND (b2103 AND (b2104 AND (b2105 AND (b2106 AND (b2107 AND (b2108 AND (b2109 AND (b2110 AND b2111))))))))))))))))))))))))))))))));
    null;
    null;
    r2114 := "0";
    null;
    r2115 := (r2114);
    r2116 := "0";
    null;
    r2117 := (r2116);
    r2118 := "0";
    null;
    r2119 := (r2118);
    r2120 := "0";
    null;
    r2121 := (r2120);
    r2122 := "0";
    null;
    r2123 := (r2122);
    r2124 := "0";
    null;
    r2125 := (r2124);
    r2126 := "0";
    null;
    r2127 := (r2126);
    r2128 := "0";
    null;
    r2129 := (r2128);
    r2130 := "0";
    null;
    r2131 := (r2130);
    r2132 := "0";
    null;
    r2133 := (r2132);
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    r2113 := (r2115 & r2117 & r2119 & r2121 & r2123 & r2125 & r2127 & r2129 & r2131 & r2133 & r2048 & r2049 & r2050 & r2051 & r2052 & r2053 & r2054 & r2055 & r2056 & r2057 & r2058 & r2059 & r2060 & r2061 & r2062 & r2063 & r2064 & r2065 & r2066 & r2067 & r2068 & r2069);
    r2046 := r2113;
    return r2046;
  end rewire_RWPreludeshiftR10_2044;
  function rewire_RWPreluderotateR19_1972(r1973 : std_logic_vector) return std_logic_vector
  is
    variable r2041 : std_logic_vector(0 to 31) := (others => '0');
    variable b2040 : boolean := false;
    variable b2039 : boolean := false;
    variable b2038 : boolean := false;
    variable b2037 : boolean := false;
    variable b2036 : boolean := false;
    variable b2035 : boolean := false;
    variable b2034 : boolean := false;
    variable b2033 : boolean := false;
    variable b2032 : boolean := false;
    variable b2031 : boolean := false;
    variable b2030 : boolean := false;
    variable b2029 : boolean := false;
    variable b2028 : boolean := false;
    variable b2027 : boolean := false;
    variable b2026 : boolean := false;
    variable b2025 : boolean := false;
    variable b2024 : boolean := false;
    variable b2023 : boolean := false;
    variable b2022 : boolean := false;
    variable b2021 : boolean := false;
    variable b2020 : boolean := false;
    variable b2019 : boolean := false;
    variable b2018 : boolean := false;
    variable b2017 : boolean := false;
    variable b2016 : boolean := false;
    variable b2015 : boolean := false;
    variable b2014 : boolean := false;
    variable b2013 : boolean := false;
    variable b2012 : boolean := false;
    variable b2011 : boolean := false;
    variable b2010 : boolean := false;
    variable b2009 : boolean := false;
    variable b2008 : boolean := false;
    variable r2007 : std_logic_vector(0 to 0) := (others => '0');
    variable r2006 : std_logic_vector(0 to 0) := (others => '0');
    variable r2005 : std_logic_vector(0 to 0) := (others => '0');
    variable r2004 : std_logic_vector(0 to 0) := (others => '0');
    variable r2003 : std_logic_vector(0 to 0) := (others => '0');
    variable r2002 : std_logic_vector(0 to 0) := (others => '0');
    variable r2001 : std_logic_vector(0 to 0) := (others => '0');
    variable r2000 : std_logic_vector(0 to 0) := (others => '0');
    variable r1999 : std_logic_vector(0 to 0) := (others => '0');
    variable r1998 : std_logic_vector(0 to 0) := (others => '0');
    variable r1997 : std_logic_vector(0 to 0) := (others => '0');
    variable r1996 : std_logic_vector(0 to 0) := (others => '0');
    variable r1995 : std_logic_vector(0 to 0) := (others => '0');
    variable r1994 : std_logic_vector(0 to 0) := (others => '0');
    variable r1993 : std_logic_vector(0 to 0) := (others => '0');
    variable r1992 : std_logic_vector(0 to 0) := (others => '0');
    variable r1991 : std_logic_vector(0 to 0) := (others => '0');
    variable r1990 : std_logic_vector(0 to 0) := (others => '0');
    variable r1989 : std_logic_vector(0 to 0) := (others => '0');
    variable r1988 : std_logic_vector(0 to 0) := (others => '0');
    variable r1987 : std_logic_vector(0 to 0) := (others => '0');
    variable r1986 : std_logic_vector(0 to 0) := (others => '0');
    variable r1985 : std_logic_vector(0 to 0) := (others => '0');
    variable r1984 : std_logic_vector(0 to 0) := (others => '0');
    variable r1983 : std_logic_vector(0 to 0) := (others => '0');
    variable r1982 : std_logic_vector(0 to 0) := (others => '0');
    variable r1981 : std_logic_vector(0 to 0) := (others => '0');
    variable r1980 : std_logic_vector(0 to 0) := (others => '0');
    variable r1979 : std_logic_vector(0 to 0) := (others => '0');
    variable r1978 : std_logic_vector(0 to 0) := (others => '0');
    variable r1977 : std_logic_vector(0 to 0) := (others => '0');
    variable r1976 : std_logic_vector(0 to 0) := (others => '0');
    variable b1975 : boolean := false;
    variable r1974 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    b1975 := true;
    r1976 := r1973(0 to 0);
    r1977 := r1973(1 to 1);
    r1978 := r1973(2 to 2);
    r1979 := r1973(3 to 3);
    r1980 := r1973(4 to 4);
    r1981 := r1973(5 to 5);
    r1982 := r1973(6 to 6);
    r1983 := r1973(7 to 7);
    r1984 := r1973(8 to 8);
    r1985 := r1973(9 to 9);
    r1986 := r1973(10 to 10);
    r1987 := r1973(11 to 11);
    r1988 := r1973(12 to 12);
    r1989 := r1973(13 to 13);
    r1990 := r1973(14 to 14);
    r1991 := r1973(15 to 15);
    r1992 := r1973(16 to 16);
    r1993 := r1973(17 to 17);
    r1994 := r1973(18 to 18);
    r1995 := r1973(19 to 19);
    r1996 := r1973(20 to 20);
    r1997 := r1973(21 to 21);
    r1998 := r1973(22 to 22);
    r1999 := r1973(23 to 23);
    r2000 := r1973(24 to 24);
    r2001 := r1973(25 to 25);
    r2002 := r1973(26 to 26);
    r2003 := r1973(27 to 27);
    r2004 := r1973(28 to 28);
    r2005 := r1973(29 to 29);
    r2006 := r1973(30 to 30);
    r2007 := r1973(31 to 31);
    b2008 := true;
    b2009 := true;
    b2010 := true;
    b2011 := true;
    b2012 := true;
    b2013 := true;
    b2014 := true;
    b2015 := true;
    b2016 := true;
    b2017 := true;
    b2018 := true;
    b2019 := true;
    b2020 := true;
    b2021 := true;
    b2022 := true;
    b2023 := true;
    b2024 := true;
    b2025 := true;
    b2026 := true;
    b2027 := true;
    b2028 := true;
    b2029 := true;
    b2030 := true;
    b2031 := true;
    b2032 := true;
    b2033 := true;
    b2034 := true;
    b2035 := true;
    b2036 := true;
    b2037 := true;
    b2038 := true;
    b2039 := true;
    b2040 := (b1975 AND (b2008 AND (b2009 AND (b2010 AND (b2011 AND (b2012 AND (b2013 AND (b2014 AND (b2015 AND (b2016 AND (b2017 AND (b2018 AND (b2019 AND (b2020 AND (b2021 AND (b2022 AND (b2023 AND (b2024 AND (b2025 AND (b2026 AND (b2027 AND (b2028 AND (b2029 AND (b2030 AND (b2031 AND (b2032 AND (b2033 AND (b2034 AND (b2035 AND (b2036 AND (b2037 AND (b2038 AND b2039))))))))))))))))))))))))))))))));
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    r2041 := (r1989 & r1990 & r1991 & r1992 & r1993 & r1994 & r1995 & r1996 & r1997 & r1998 & r1999 & r2000 & r2001 & r2002 & r2003 & r2004 & r2005 & r2006 & r2007 & r1976 & r1977 & r1978 & r1979 & r1980 & r1981 & r1982 & r1983 & r1984 & r1985 & r1986 & r1987 & r1988);
    r1974 := r2041;
    return r1974;
  end rewire_RWPreluderotateR19_1972;
  function rewire_RWPreluderotateR17_1901(r1902 : std_logic_vector) return std_logic_vector
  is
    variable r1970 : std_logic_vector(0 to 31) := (others => '0');
    variable b1969 : boolean := false;
    variable b1968 : boolean := false;
    variable b1967 : boolean := false;
    variable b1966 : boolean := false;
    variable b1965 : boolean := false;
    variable b1964 : boolean := false;
    variable b1963 : boolean := false;
    variable b1962 : boolean := false;
    variable b1961 : boolean := false;
    variable b1960 : boolean := false;
    variable b1959 : boolean := false;
    variable b1958 : boolean := false;
    variable b1957 : boolean := false;
    variable b1956 : boolean := false;
    variable b1955 : boolean := false;
    variable b1954 : boolean := false;
    variable b1953 : boolean := false;
    variable b1952 : boolean := false;
    variable b1951 : boolean := false;
    variable b1950 : boolean := false;
    variable b1949 : boolean := false;
    variable b1948 : boolean := false;
    variable b1947 : boolean := false;
    variable b1946 : boolean := false;
    variable b1945 : boolean := false;
    variable b1944 : boolean := false;
    variable b1943 : boolean := false;
    variable b1942 : boolean := false;
    variable b1941 : boolean := false;
    variable b1940 : boolean := false;
    variable b1939 : boolean := false;
    variable b1938 : boolean := false;
    variable b1937 : boolean := false;
    variable r1936 : std_logic_vector(0 to 0) := (others => '0');
    variable r1935 : std_logic_vector(0 to 0) := (others => '0');
    variable r1934 : std_logic_vector(0 to 0) := (others => '0');
    variable r1933 : std_logic_vector(0 to 0) := (others => '0');
    variable r1932 : std_logic_vector(0 to 0) := (others => '0');
    variable r1931 : std_logic_vector(0 to 0) := (others => '0');
    variable r1930 : std_logic_vector(0 to 0) := (others => '0');
    variable r1929 : std_logic_vector(0 to 0) := (others => '0');
    variable r1928 : std_logic_vector(0 to 0) := (others => '0');
    variable r1927 : std_logic_vector(0 to 0) := (others => '0');
    variable r1926 : std_logic_vector(0 to 0) := (others => '0');
    variable r1925 : std_logic_vector(0 to 0) := (others => '0');
    variable r1924 : std_logic_vector(0 to 0) := (others => '0');
    variable r1923 : std_logic_vector(0 to 0) := (others => '0');
    variable r1922 : std_logic_vector(0 to 0) := (others => '0');
    variable r1921 : std_logic_vector(0 to 0) := (others => '0');
    variable r1920 : std_logic_vector(0 to 0) := (others => '0');
    variable r1919 : std_logic_vector(0 to 0) := (others => '0');
    variable r1918 : std_logic_vector(0 to 0) := (others => '0');
    variable r1917 : std_logic_vector(0 to 0) := (others => '0');
    variable r1916 : std_logic_vector(0 to 0) := (others => '0');
    variable r1915 : std_logic_vector(0 to 0) := (others => '0');
    variable r1914 : std_logic_vector(0 to 0) := (others => '0');
    variable r1913 : std_logic_vector(0 to 0) := (others => '0');
    variable r1912 : std_logic_vector(0 to 0) := (others => '0');
    variable r1911 : std_logic_vector(0 to 0) := (others => '0');
    variable r1910 : std_logic_vector(0 to 0) := (others => '0');
    variable r1909 : std_logic_vector(0 to 0) := (others => '0');
    variable r1908 : std_logic_vector(0 to 0) := (others => '0');
    variable r1907 : std_logic_vector(0 to 0) := (others => '0');
    variable r1906 : std_logic_vector(0 to 0) := (others => '0');
    variable r1905 : std_logic_vector(0 to 0) := (others => '0');
    variable b1904 : boolean := false;
    variable r1903 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    b1904 := true;
    r1905 := r1902(0 to 0);
    r1906 := r1902(1 to 1);
    r1907 := r1902(2 to 2);
    r1908 := r1902(3 to 3);
    r1909 := r1902(4 to 4);
    r1910 := r1902(5 to 5);
    r1911 := r1902(6 to 6);
    r1912 := r1902(7 to 7);
    r1913 := r1902(8 to 8);
    r1914 := r1902(9 to 9);
    r1915 := r1902(10 to 10);
    r1916 := r1902(11 to 11);
    r1917 := r1902(12 to 12);
    r1918 := r1902(13 to 13);
    r1919 := r1902(14 to 14);
    r1920 := r1902(15 to 15);
    r1921 := r1902(16 to 16);
    r1922 := r1902(17 to 17);
    r1923 := r1902(18 to 18);
    r1924 := r1902(19 to 19);
    r1925 := r1902(20 to 20);
    r1926 := r1902(21 to 21);
    r1927 := r1902(22 to 22);
    r1928 := r1902(23 to 23);
    r1929 := r1902(24 to 24);
    r1930 := r1902(25 to 25);
    r1931 := r1902(26 to 26);
    r1932 := r1902(27 to 27);
    r1933 := r1902(28 to 28);
    r1934 := r1902(29 to 29);
    r1935 := r1902(30 to 30);
    r1936 := r1902(31 to 31);
    b1937 := true;
    b1938 := true;
    b1939 := true;
    b1940 := true;
    b1941 := true;
    b1942 := true;
    b1943 := true;
    b1944 := true;
    b1945 := true;
    b1946 := true;
    b1947 := true;
    b1948 := true;
    b1949 := true;
    b1950 := true;
    b1951 := true;
    b1952 := true;
    b1953 := true;
    b1954 := true;
    b1955 := true;
    b1956 := true;
    b1957 := true;
    b1958 := true;
    b1959 := true;
    b1960 := true;
    b1961 := true;
    b1962 := true;
    b1963 := true;
    b1964 := true;
    b1965 := true;
    b1966 := true;
    b1967 := true;
    b1968 := true;
    b1969 := (b1904 AND (b1937 AND (b1938 AND (b1939 AND (b1940 AND (b1941 AND (b1942 AND (b1943 AND (b1944 AND (b1945 AND (b1946 AND (b1947 AND (b1948 AND (b1949 AND (b1950 AND (b1951 AND (b1952 AND (b1953 AND (b1954 AND (b1955 AND (b1956 AND (b1957 AND (b1958 AND (b1959 AND (b1960 AND (b1961 AND (b1962 AND (b1963 AND (b1964 AND (b1965 AND (b1966 AND (b1967 AND b1968))))))))))))))))))))))))))))))));
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    r1970 := (r1920 & r1921 & r1922 & r1923 & r1924 & r1925 & r1926 & r1927 & r1928 & r1929 & r1930 & r1931 & r1932 & r1933 & r1934 & r1935 & r1936 & r1905 & r1906 & r1907 & r1908 & r1909 & r1910 & r1911 & r1912 & r1913 & r1914 & r1915 & r1916 & r1917 & r1918 & r1919);
    r1903 := r1970;
    return r1903;
  end rewire_RWPreluderotateR17_1901;
  function rewire_MaininitialSHA256State_28 return std_logic_vector
  is
    variable r565 : std_logic_vector(0 to 31) := (others => '0');
    variable r498 : std_logic_vector(0 to 31) := (others => '0');
    variable r431 : std_logic_vector(0 to 31) := (others => '0');
    variable r364 : std_logic_vector(0 to 31) := (others => '0');
    variable r297 : std_logic_vector(0 to 31) := (others => '0');
    variable r230 : std_logic_vector(0 to 31) := (others => '0');
    variable r163 : std_logic_vector(0 to 31) := (others => '0');
    variable r96 : std_logic_vector(0 to 31) := (others => '0');
    variable r29 : std_logic_vector(0 to 255) := (others => '0');
  begin
    null;
    null;
    r96 := rewire_MetaprogrammingRWw6a09e667_30;
    r163 := rewire_MetaprogrammingRWwbb67ae85_97;
    r230 := rewire_MetaprogrammingRWw3c6ef372_164;
    r297 := rewire_MetaprogrammingRWwa54ff53a_231;
    r364 := rewire_MetaprogrammingRWw510e527f_298;
    r431 := rewire_MetaprogrammingRWw9b05688c_365;
    r498 := rewire_MetaprogrammingRWw1f83d9ab_432;
    r565 := rewire_MetaprogrammingRWw5be0cd19_499;
    r29 := (r96 & r163 & r230 & r297 & r364 & r431 & r498 & r565);
    return r29;
  end rewire_MaininitialSHA256State_28;
  function rewire_MetaprogrammingRWw5be0cd19_499 return std_logic_vector
  is
    variable r564 : std_logic_vector(0 to 0) := (others => '0');
    variable r563 : std_logic_vector(0 to 0) := (others => '0');
    variable r562 : std_logic_vector(0 to 0) := (others => '0');
    variable r561 : std_logic_vector(0 to 0) := (others => '0');
    variable r560 : std_logic_vector(0 to 0) := (others => '0');
    variable r559 : std_logic_vector(0 to 0) := (others => '0');
    variable r558 : std_logic_vector(0 to 0) := (others => '0');
    variable r557 : std_logic_vector(0 to 0) := (others => '0');
    variable r556 : std_logic_vector(0 to 0) := (others => '0');
    variable r555 : std_logic_vector(0 to 0) := (others => '0');
    variable r554 : std_logic_vector(0 to 0) := (others => '0');
    variable r553 : std_logic_vector(0 to 0) := (others => '0');
    variable r552 : std_logic_vector(0 to 0) := (others => '0');
    variable r551 : std_logic_vector(0 to 0) := (others => '0');
    variable r550 : std_logic_vector(0 to 0) := (others => '0');
    variable r549 : std_logic_vector(0 to 0) := (others => '0');
    variable r548 : std_logic_vector(0 to 0) := (others => '0');
    variable r547 : std_logic_vector(0 to 0) := (others => '0');
    variable r546 : std_logic_vector(0 to 0) := (others => '0');
    variable r545 : std_logic_vector(0 to 0) := (others => '0');
    variable r544 : std_logic_vector(0 to 0) := (others => '0');
    variable r543 : std_logic_vector(0 to 0) := (others => '0');
    variable r542 : std_logic_vector(0 to 0) := (others => '0');
    variable r541 : std_logic_vector(0 to 0) := (others => '0');
    variable r540 : std_logic_vector(0 to 0) := (others => '0');
    variable r539 : std_logic_vector(0 to 0) := (others => '0');
    variable r538 : std_logic_vector(0 to 0) := (others => '0');
    variable r537 : std_logic_vector(0 to 0) := (others => '0');
    variable r536 : std_logic_vector(0 to 0) := (others => '0');
    variable r535 : std_logic_vector(0 to 0) := (others => '0');
    variable r534 : std_logic_vector(0 to 0) := (others => '0');
    variable r533 : std_logic_vector(0 to 0) := (others => '0');
    variable r532 : std_logic_vector(0 to 0) := (others => '0');
    variable r531 : std_logic_vector(0 to 0) := (others => '0');
    variable r530 : std_logic_vector(0 to 0) := (others => '0');
    variable r529 : std_logic_vector(0 to 0) := (others => '0');
    variable r528 : std_logic_vector(0 to 0) := (others => '0');
    variable r527 : std_logic_vector(0 to 0) := (others => '0');
    variable r526 : std_logic_vector(0 to 0) := (others => '0');
    variable r525 : std_logic_vector(0 to 0) := (others => '0');
    variable r524 : std_logic_vector(0 to 0) := (others => '0');
    variable r523 : std_logic_vector(0 to 0) := (others => '0');
    variable r522 : std_logic_vector(0 to 0) := (others => '0');
    variable r521 : std_logic_vector(0 to 0) := (others => '0');
    variable r520 : std_logic_vector(0 to 0) := (others => '0');
    variable r519 : std_logic_vector(0 to 0) := (others => '0');
    variable r518 : std_logic_vector(0 to 0) := (others => '0');
    variable r517 : std_logic_vector(0 to 0) := (others => '0');
    variable r516 : std_logic_vector(0 to 0) := (others => '0');
    variable r515 : std_logic_vector(0 to 0) := (others => '0');
    variable r514 : std_logic_vector(0 to 0) := (others => '0');
    variable r513 : std_logic_vector(0 to 0) := (others => '0');
    variable r512 : std_logic_vector(0 to 0) := (others => '0');
    variable r511 : std_logic_vector(0 to 0) := (others => '0');
    variable r510 : std_logic_vector(0 to 0) := (others => '0');
    variable r509 : std_logic_vector(0 to 0) := (others => '0');
    variable r508 : std_logic_vector(0 to 0) := (others => '0');
    variable r507 : std_logic_vector(0 to 0) := (others => '0');
    variable r506 : std_logic_vector(0 to 0) := (others => '0');
    variable r505 : std_logic_vector(0 to 0) := (others => '0');
    variable r504 : std_logic_vector(0 to 0) := (others => '0');
    variable r503 : std_logic_vector(0 to 0) := (others => '0');
    variable r502 : std_logic_vector(0 to 0) := (others => '0');
    variable r501 : std_logic_vector(0 to 0) := (others => '0');
    variable r500 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r501 := "0";
    null;
    r502 := (r501);
    r503 := "1";
    null;
    r504 := (r503);
    r505 := "0";
    null;
    r506 := (r505);
    r507 := "1";
    null;
    r508 := (r507);
    r509 := "1";
    null;
    r510 := (r509);
    r511 := "0";
    null;
    r512 := (r511);
    r513 := "1";
    null;
    r514 := (r513);
    r515 := "1";
    null;
    r516 := (r515);
    r517 := "1";
    null;
    r518 := (r517);
    r519 := "1";
    null;
    r520 := (r519);
    r521 := "1";
    null;
    r522 := (r521);
    r523 := "0";
    null;
    r524 := (r523);
    r525 := "0";
    null;
    r526 := (r525);
    r527 := "0";
    null;
    r528 := (r527);
    r529 := "0";
    null;
    r530 := (r529);
    r531 := "0";
    null;
    r532 := (r531);
    r533 := "1";
    null;
    r534 := (r533);
    r535 := "1";
    null;
    r536 := (r535);
    r537 := "0";
    null;
    r538 := (r537);
    r539 := "0";
    null;
    r540 := (r539);
    r541 := "1";
    null;
    r542 := (r541);
    r543 := "1";
    null;
    r544 := (r543);
    r545 := "0";
    null;
    r546 := (r545);
    r547 := "1";
    null;
    r548 := (r547);
    r549 := "0";
    null;
    r550 := (r549);
    r551 := "0";
    null;
    r552 := (r551);
    r553 := "0";
    null;
    r554 := (r553);
    r555 := "1";
    null;
    r556 := (r555);
    r557 := "1";
    null;
    r558 := (r557);
    r559 := "0";
    null;
    r560 := (r559);
    r561 := "0";
    null;
    r562 := (r561);
    r563 := "1";
    null;
    r564 := (r563);
    r500 := (r502 & r504 & r506 & r508 & r510 & r512 & r514 & r516 & r518 & r520 & r522 & r524 & r526 & r528 & r530 & r532 & r534 & r536 & r538 & r540 & r542 & r544 & r546 & r548 & r550 & r552 & r554 & r556 & r558 & r560 & r562 & r564);
    return r500;
  end rewire_MetaprogrammingRWw5be0cd19_499;
  function rewire_MetaprogrammingRWw1f83d9ab_432 return std_logic_vector
  is
    variable r497 : std_logic_vector(0 to 0) := (others => '0');
    variable r496 : std_logic_vector(0 to 0) := (others => '0');
    variable r495 : std_logic_vector(0 to 0) := (others => '0');
    variable r494 : std_logic_vector(0 to 0) := (others => '0');
    variable r493 : std_logic_vector(0 to 0) := (others => '0');
    variable r492 : std_logic_vector(0 to 0) := (others => '0');
    variable r491 : std_logic_vector(0 to 0) := (others => '0');
    variable r490 : std_logic_vector(0 to 0) := (others => '0');
    variable r489 : std_logic_vector(0 to 0) := (others => '0');
    variable r488 : std_logic_vector(0 to 0) := (others => '0');
    variable r487 : std_logic_vector(0 to 0) := (others => '0');
    variable r486 : std_logic_vector(0 to 0) := (others => '0');
    variable r485 : std_logic_vector(0 to 0) := (others => '0');
    variable r484 : std_logic_vector(0 to 0) := (others => '0');
    variable r483 : std_logic_vector(0 to 0) := (others => '0');
    variable r482 : std_logic_vector(0 to 0) := (others => '0');
    variable r481 : std_logic_vector(0 to 0) := (others => '0');
    variable r480 : std_logic_vector(0 to 0) := (others => '0');
    variable r479 : std_logic_vector(0 to 0) := (others => '0');
    variable r478 : std_logic_vector(0 to 0) := (others => '0');
    variable r477 : std_logic_vector(0 to 0) := (others => '0');
    variable r476 : std_logic_vector(0 to 0) := (others => '0');
    variable r475 : std_logic_vector(0 to 0) := (others => '0');
    variable r474 : std_logic_vector(0 to 0) := (others => '0');
    variable r473 : std_logic_vector(0 to 0) := (others => '0');
    variable r472 : std_logic_vector(0 to 0) := (others => '0');
    variable r471 : std_logic_vector(0 to 0) := (others => '0');
    variable r470 : std_logic_vector(0 to 0) := (others => '0');
    variable r469 : std_logic_vector(0 to 0) := (others => '0');
    variable r468 : std_logic_vector(0 to 0) := (others => '0');
    variable r467 : std_logic_vector(0 to 0) := (others => '0');
    variable r466 : std_logic_vector(0 to 0) := (others => '0');
    variable r465 : std_logic_vector(0 to 0) := (others => '0');
    variable r464 : std_logic_vector(0 to 0) := (others => '0');
    variable r463 : std_logic_vector(0 to 0) := (others => '0');
    variable r462 : std_logic_vector(0 to 0) := (others => '0');
    variable r461 : std_logic_vector(0 to 0) := (others => '0');
    variable r460 : std_logic_vector(0 to 0) := (others => '0');
    variable r459 : std_logic_vector(0 to 0) := (others => '0');
    variable r458 : std_logic_vector(0 to 0) := (others => '0');
    variable r457 : std_logic_vector(0 to 0) := (others => '0');
    variable r456 : std_logic_vector(0 to 0) := (others => '0');
    variable r455 : std_logic_vector(0 to 0) := (others => '0');
    variable r454 : std_logic_vector(0 to 0) := (others => '0');
    variable r453 : std_logic_vector(0 to 0) := (others => '0');
    variable r452 : std_logic_vector(0 to 0) := (others => '0');
    variable r451 : std_logic_vector(0 to 0) := (others => '0');
    variable r450 : std_logic_vector(0 to 0) := (others => '0');
    variable r449 : std_logic_vector(0 to 0) := (others => '0');
    variable r448 : std_logic_vector(0 to 0) := (others => '0');
    variable r447 : std_logic_vector(0 to 0) := (others => '0');
    variable r446 : std_logic_vector(0 to 0) := (others => '0');
    variable r445 : std_logic_vector(0 to 0) := (others => '0');
    variable r444 : std_logic_vector(0 to 0) := (others => '0');
    variable r443 : std_logic_vector(0 to 0) := (others => '0');
    variable r442 : std_logic_vector(0 to 0) := (others => '0');
    variable r441 : std_logic_vector(0 to 0) := (others => '0');
    variable r440 : std_logic_vector(0 to 0) := (others => '0');
    variable r439 : std_logic_vector(0 to 0) := (others => '0');
    variable r438 : std_logic_vector(0 to 0) := (others => '0');
    variable r437 : std_logic_vector(0 to 0) := (others => '0');
    variable r436 : std_logic_vector(0 to 0) := (others => '0');
    variable r435 : std_logic_vector(0 to 0) := (others => '0');
    variable r434 : std_logic_vector(0 to 0) := (others => '0');
    variable r433 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r434 := "0";
    null;
    r435 := (r434);
    r436 := "0";
    null;
    r437 := (r436);
    r438 := "0";
    null;
    r439 := (r438);
    r440 := "1";
    null;
    r441 := (r440);
    r442 := "1";
    null;
    r443 := (r442);
    r444 := "1";
    null;
    r445 := (r444);
    r446 := "1";
    null;
    r447 := (r446);
    r448 := "1";
    null;
    r449 := (r448);
    r450 := "1";
    null;
    r451 := (r450);
    r452 := "0";
    null;
    r453 := (r452);
    r454 := "0";
    null;
    r455 := (r454);
    r456 := "0";
    null;
    r457 := (r456);
    r458 := "0";
    null;
    r459 := (r458);
    r460 := "0";
    null;
    r461 := (r460);
    r462 := "1";
    null;
    r463 := (r462);
    r464 := "1";
    null;
    r465 := (r464);
    r466 := "1";
    null;
    r467 := (r466);
    r468 := "1";
    null;
    r469 := (r468);
    r470 := "0";
    null;
    r471 := (r470);
    r472 := "1";
    null;
    r473 := (r472);
    r474 := "1";
    null;
    r475 := (r474);
    r476 := "0";
    null;
    r477 := (r476);
    r478 := "0";
    null;
    r479 := (r478);
    r480 := "1";
    null;
    r481 := (r480);
    r482 := "1";
    null;
    r483 := (r482);
    r484 := "0";
    null;
    r485 := (r484);
    r486 := "1";
    null;
    r487 := (r486);
    r488 := "0";
    null;
    r489 := (r488);
    r490 := "1";
    null;
    r491 := (r490);
    r492 := "0";
    null;
    r493 := (r492);
    r494 := "1";
    null;
    r495 := (r494);
    r496 := "1";
    null;
    r497 := (r496);
    r433 := (r435 & r437 & r439 & r441 & r443 & r445 & r447 & r449 & r451 & r453 & r455 & r457 & r459 & r461 & r463 & r465 & r467 & r469 & r471 & r473 & r475 & r477 & r479 & r481 & r483 & r485 & r487 & r489 & r491 & r493 & r495 & r497);
    return r433;
  end rewire_MetaprogrammingRWw1f83d9ab_432;
  function rewire_MetaprogrammingRWw9b05688c_365 return std_logic_vector
  is
    variable r430 : std_logic_vector(0 to 0) := (others => '0');
    variable r429 : std_logic_vector(0 to 0) := (others => '0');
    variable r428 : std_logic_vector(0 to 0) := (others => '0');
    variable r427 : std_logic_vector(0 to 0) := (others => '0');
    variable r426 : std_logic_vector(0 to 0) := (others => '0');
    variable r425 : std_logic_vector(0 to 0) := (others => '0');
    variable r424 : std_logic_vector(0 to 0) := (others => '0');
    variable r423 : std_logic_vector(0 to 0) := (others => '0');
    variable r422 : std_logic_vector(0 to 0) := (others => '0');
    variable r421 : std_logic_vector(0 to 0) := (others => '0');
    variable r420 : std_logic_vector(0 to 0) := (others => '0');
    variable r419 : std_logic_vector(0 to 0) := (others => '0');
    variable r418 : std_logic_vector(0 to 0) := (others => '0');
    variable r417 : std_logic_vector(0 to 0) := (others => '0');
    variable r416 : std_logic_vector(0 to 0) := (others => '0');
    variable r415 : std_logic_vector(0 to 0) := (others => '0');
    variable r414 : std_logic_vector(0 to 0) := (others => '0');
    variable r413 : std_logic_vector(0 to 0) := (others => '0');
    variable r412 : std_logic_vector(0 to 0) := (others => '0');
    variable r411 : std_logic_vector(0 to 0) := (others => '0');
    variable r410 : std_logic_vector(0 to 0) := (others => '0');
    variable r409 : std_logic_vector(0 to 0) := (others => '0');
    variable r408 : std_logic_vector(0 to 0) := (others => '0');
    variable r407 : std_logic_vector(0 to 0) := (others => '0');
    variable r406 : std_logic_vector(0 to 0) := (others => '0');
    variable r405 : std_logic_vector(0 to 0) := (others => '0');
    variable r404 : std_logic_vector(0 to 0) := (others => '0');
    variable r403 : std_logic_vector(0 to 0) := (others => '0');
    variable r402 : std_logic_vector(0 to 0) := (others => '0');
    variable r401 : std_logic_vector(0 to 0) := (others => '0');
    variable r400 : std_logic_vector(0 to 0) := (others => '0');
    variable r399 : std_logic_vector(0 to 0) := (others => '0');
    variable r398 : std_logic_vector(0 to 0) := (others => '0');
    variable r397 : std_logic_vector(0 to 0) := (others => '0');
    variable r396 : std_logic_vector(0 to 0) := (others => '0');
    variable r395 : std_logic_vector(0 to 0) := (others => '0');
    variable r394 : std_logic_vector(0 to 0) := (others => '0');
    variable r393 : std_logic_vector(0 to 0) := (others => '0');
    variable r392 : std_logic_vector(0 to 0) := (others => '0');
    variable r391 : std_logic_vector(0 to 0) := (others => '0');
    variable r390 : std_logic_vector(0 to 0) := (others => '0');
    variable r389 : std_logic_vector(0 to 0) := (others => '0');
    variable r388 : std_logic_vector(0 to 0) := (others => '0');
    variable r387 : std_logic_vector(0 to 0) := (others => '0');
    variable r386 : std_logic_vector(0 to 0) := (others => '0');
    variable r385 : std_logic_vector(0 to 0) := (others => '0');
    variable r384 : std_logic_vector(0 to 0) := (others => '0');
    variable r383 : std_logic_vector(0 to 0) := (others => '0');
    variable r382 : std_logic_vector(0 to 0) := (others => '0');
    variable r381 : std_logic_vector(0 to 0) := (others => '0');
    variable r380 : std_logic_vector(0 to 0) := (others => '0');
    variable r379 : std_logic_vector(0 to 0) := (others => '0');
    variable r378 : std_logic_vector(0 to 0) := (others => '0');
    variable r377 : std_logic_vector(0 to 0) := (others => '0');
    variable r376 : std_logic_vector(0 to 0) := (others => '0');
    variable r375 : std_logic_vector(0 to 0) := (others => '0');
    variable r374 : std_logic_vector(0 to 0) := (others => '0');
    variable r373 : std_logic_vector(0 to 0) := (others => '0');
    variable r372 : std_logic_vector(0 to 0) := (others => '0');
    variable r371 : std_logic_vector(0 to 0) := (others => '0');
    variable r370 : std_logic_vector(0 to 0) := (others => '0');
    variable r369 : std_logic_vector(0 to 0) := (others => '0');
    variable r368 : std_logic_vector(0 to 0) := (others => '0');
    variable r367 : std_logic_vector(0 to 0) := (others => '0');
    variable r366 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r367 := "1";
    null;
    r368 := (r367);
    r369 := "0";
    null;
    r370 := (r369);
    r371 := "0";
    null;
    r372 := (r371);
    r373 := "1";
    null;
    r374 := (r373);
    r375 := "1";
    null;
    r376 := (r375);
    r377 := "0";
    null;
    r378 := (r377);
    r379 := "1";
    null;
    r380 := (r379);
    r381 := "1";
    null;
    r382 := (r381);
    r383 := "0";
    null;
    r384 := (r383);
    r385 := "0";
    null;
    r386 := (r385);
    r387 := "0";
    null;
    r388 := (r387);
    r389 := "0";
    null;
    r390 := (r389);
    r391 := "0";
    null;
    r392 := (r391);
    r393 := "1";
    null;
    r394 := (r393);
    r395 := "0";
    null;
    r396 := (r395);
    r397 := "1";
    null;
    r398 := (r397);
    r399 := "0";
    null;
    r400 := (r399);
    r401 := "1";
    null;
    r402 := (r401);
    r403 := "1";
    null;
    r404 := (r403);
    r405 := "0";
    null;
    r406 := (r405);
    r407 := "1";
    null;
    r408 := (r407);
    r409 := "0";
    null;
    r410 := (r409);
    r411 := "0";
    null;
    r412 := (r411);
    r413 := "0";
    null;
    r414 := (r413);
    r415 := "1";
    null;
    r416 := (r415);
    r417 := "0";
    null;
    r418 := (r417);
    r419 := "0";
    null;
    r420 := (r419);
    r421 := "0";
    null;
    r422 := (r421);
    r423 := "1";
    null;
    r424 := (r423);
    r425 := "1";
    null;
    r426 := (r425);
    r427 := "0";
    null;
    r428 := (r427);
    r429 := "0";
    null;
    r430 := (r429);
    r366 := (r368 & r370 & r372 & r374 & r376 & r378 & r380 & r382 & r384 & r386 & r388 & r390 & r392 & r394 & r396 & r398 & r400 & r402 & r404 & r406 & r408 & r410 & r412 & r414 & r416 & r418 & r420 & r422 & r424 & r426 & r428 & r430);
    return r366;
  end rewire_MetaprogrammingRWw9b05688c_365;
  function rewire_MetaprogrammingRWw510e527f_298 return std_logic_vector
  is
    variable r363 : std_logic_vector(0 to 0) := (others => '0');
    variable r362 : std_logic_vector(0 to 0) := (others => '0');
    variable r361 : std_logic_vector(0 to 0) := (others => '0');
    variable r360 : std_logic_vector(0 to 0) := (others => '0');
    variable r359 : std_logic_vector(0 to 0) := (others => '0');
    variable r358 : std_logic_vector(0 to 0) := (others => '0');
    variable r357 : std_logic_vector(0 to 0) := (others => '0');
    variable r356 : std_logic_vector(0 to 0) := (others => '0');
    variable r355 : std_logic_vector(0 to 0) := (others => '0');
    variable r354 : std_logic_vector(0 to 0) := (others => '0');
    variable r353 : std_logic_vector(0 to 0) := (others => '0');
    variable r352 : std_logic_vector(0 to 0) := (others => '0');
    variable r351 : std_logic_vector(0 to 0) := (others => '0');
    variable r350 : std_logic_vector(0 to 0) := (others => '0');
    variable r349 : std_logic_vector(0 to 0) := (others => '0');
    variable r348 : std_logic_vector(0 to 0) := (others => '0');
    variable r347 : std_logic_vector(0 to 0) := (others => '0');
    variable r346 : std_logic_vector(0 to 0) := (others => '0');
    variable r345 : std_logic_vector(0 to 0) := (others => '0');
    variable r344 : std_logic_vector(0 to 0) := (others => '0');
    variable r343 : std_logic_vector(0 to 0) := (others => '0');
    variable r342 : std_logic_vector(0 to 0) := (others => '0');
    variable r341 : std_logic_vector(0 to 0) := (others => '0');
    variable r340 : std_logic_vector(0 to 0) := (others => '0');
    variable r339 : std_logic_vector(0 to 0) := (others => '0');
    variable r338 : std_logic_vector(0 to 0) := (others => '0');
    variable r337 : std_logic_vector(0 to 0) := (others => '0');
    variable r336 : std_logic_vector(0 to 0) := (others => '0');
    variable r335 : std_logic_vector(0 to 0) := (others => '0');
    variable r334 : std_logic_vector(0 to 0) := (others => '0');
    variable r333 : std_logic_vector(0 to 0) := (others => '0');
    variable r332 : std_logic_vector(0 to 0) := (others => '0');
    variable r331 : std_logic_vector(0 to 0) := (others => '0');
    variable r330 : std_logic_vector(0 to 0) := (others => '0');
    variable r329 : std_logic_vector(0 to 0) := (others => '0');
    variable r328 : std_logic_vector(0 to 0) := (others => '0');
    variable r327 : std_logic_vector(0 to 0) := (others => '0');
    variable r326 : std_logic_vector(0 to 0) := (others => '0');
    variable r325 : std_logic_vector(0 to 0) := (others => '0');
    variable r324 : std_logic_vector(0 to 0) := (others => '0');
    variable r323 : std_logic_vector(0 to 0) := (others => '0');
    variable r322 : std_logic_vector(0 to 0) := (others => '0');
    variable r321 : std_logic_vector(0 to 0) := (others => '0');
    variable r320 : std_logic_vector(0 to 0) := (others => '0');
    variable r319 : std_logic_vector(0 to 0) := (others => '0');
    variable r318 : std_logic_vector(0 to 0) := (others => '0');
    variable r317 : std_logic_vector(0 to 0) := (others => '0');
    variable r316 : std_logic_vector(0 to 0) := (others => '0');
    variable r315 : std_logic_vector(0 to 0) := (others => '0');
    variable r314 : std_logic_vector(0 to 0) := (others => '0');
    variable r313 : std_logic_vector(0 to 0) := (others => '0');
    variable r312 : std_logic_vector(0 to 0) := (others => '0');
    variable r311 : std_logic_vector(0 to 0) := (others => '0');
    variable r310 : std_logic_vector(0 to 0) := (others => '0');
    variable r309 : std_logic_vector(0 to 0) := (others => '0');
    variable r308 : std_logic_vector(0 to 0) := (others => '0');
    variable r307 : std_logic_vector(0 to 0) := (others => '0');
    variable r306 : std_logic_vector(0 to 0) := (others => '0');
    variable r305 : std_logic_vector(0 to 0) := (others => '0');
    variable r304 : std_logic_vector(0 to 0) := (others => '0');
    variable r303 : std_logic_vector(0 to 0) := (others => '0');
    variable r302 : std_logic_vector(0 to 0) := (others => '0');
    variable r301 : std_logic_vector(0 to 0) := (others => '0');
    variable r300 : std_logic_vector(0 to 0) := (others => '0');
    variable r299 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r300 := "0";
    null;
    r301 := (r300);
    r302 := "1";
    null;
    r303 := (r302);
    r304 := "0";
    null;
    r305 := (r304);
    r306 := "1";
    null;
    r307 := (r306);
    r308 := "0";
    null;
    r309 := (r308);
    r310 := "0";
    null;
    r311 := (r310);
    r312 := "0";
    null;
    r313 := (r312);
    r314 := "1";
    null;
    r315 := (r314);
    r316 := "0";
    null;
    r317 := (r316);
    r318 := "0";
    null;
    r319 := (r318);
    r320 := "0";
    null;
    r321 := (r320);
    r322 := "0";
    null;
    r323 := (r322);
    r324 := "1";
    null;
    r325 := (r324);
    r326 := "1";
    null;
    r327 := (r326);
    r328 := "1";
    null;
    r329 := (r328);
    r330 := "0";
    null;
    r331 := (r330);
    r332 := "0";
    null;
    r333 := (r332);
    r334 := "1";
    null;
    r335 := (r334);
    r336 := "0";
    null;
    r337 := (r336);
    r338 := "1";
    null;
    r339 := (r338);
    r340 := "0";
    null;
    r341 := (r340);
    r342 := "0";
    null;
    r343 := (r342);
    r344 := "1";
    null;
    r345 := (r344);
    r346 := "0";
    null;
    r347 := (r346);
    r348 := "0";
    null;
    r349 := (r348);
    r350 := "1";
    null;
    r351 := (r350);
    r352 := "1";
    null;
    r353 := (r352);
    r354 := "1";
    null;
    r355 := (r354);
    r356 := "1";
    null;
    r357 := (r356);
    r358 := "1";
    null;
    r359 := (r358);
    r360 := "1";
    null;
    r361 := (r360);
    r362 := "1";
    null;
    r363 := (r362);
    r299 := (r301 & r303 & r305 & r307 & r309 & r311 & r313 & r315 & r317 & r319 & r321 & r323 & r325 & r327 & r329 & r331 & r333 & r335 & r337 & r339 & r341 & r343 & r345 & r347 & r349 & r351 & r353 & r355 & r357 & r359 & r361 & r363);
    return r299;
  end rewire_MetaprogrammingRWw510e527f_298;
  function rewire_MetaprogrammingRWwa54ff53a_231 return std_logic_vector
  is
    variable r296 : std_logic_vector(0 to 0) := (others => '0');
    variable r295 : std_logic_vector(0 to 0) := (others => '0');
    variable r294 : std_logic_vector(0 to 0) := (others => '0');
    variable r293 : std_logic_vector(0 to 0) := (others => '0');
    variable r292 : std_logic_vector(0 to 0) := (others => '0');
    variable r291 : std_logic_vector(0 to 0) := (others => '0');
    variable r290 : std_logic_vector(0 to 0) := (others => '0');
    variable r289 : std_logic_vector(0 to 0) := (others => '0');
    variable r288 : std_logic_vector(0 to 0) := (others => '0');
    variable r287 : std_logic_vector(0 to 0) := (others => '0');
    variable r286 : std_logic_vector(0 to 0) := (others => '0');
    variable r285 : std_logic_vector(0 to 0) := (others => '0');
    variable r284 : std_logic_vector(0 to 0) := (others => '0');
    variable r283 : std_logic_vector(0 to 0) := (others => '0');
    variable r282 : std_logic_vector(0 to 0) := (others => '0');
    variable r281 : std_logic_vector(0 to 0) := (others => '0');
    variable r280 : std_logic_vector(0 to 0) := (others => '0');
    variable r279 : std_logic_vector(0 to 0) := (others => '0');
    variable r278 : std_logic_vector(0 to 0) := (others => '0');
    variable r277 : std_logic_vector(0 to 0) := (others => '0');
    variable r276 : std_logic_vector(0 to 0) := (others => '0');
    variable r275 : std_logic_vector(0 to 0) := (others => '0');
    variable r274 : std_logic_vector(0 to 0) := (others => '0');
    variable r273 : std_logic_vector(0 to 0) := (others => '0');
    variable r272 : std_logic_vector(0 to 0) := (others => '0');
    variable r271 : std_logic_vector(0 to 0) := (others => '0');
    variable r270 : std_logic_vector(0 to 0) := (others => '0');
    variable r269 : std_logic_vector(0 to 0) := (others => '0');
    variable r268 : std_logic_vector(0 to 0) := (others => '0');
    variable r267 : std_logic_vector(0 to 0) := (others => '0');
    variable r266 : std_logic_vector(0 to 0) := (others => '0');
    variable r265 : std_logic_vector(0 to 0) := (others => '0');
    variable r264 : std_logic_vector(0 to 0) := (others => '0');
    variable r263 : std_logic_vector(0 to 0) := (others => '0');
    variable r262 : std_logic_vector(0 to 0) := (others => '0');
    variable r261 : std_logic_vector(0 to 0) := (others => '0');
    variable r260 : std_logic_vector(0 to 0) := (others => '0');
    variable r259 : std_logic_vector(0 to 0) := (others => '0');
    variable r258 : std_logic_vector(0 to 0) := (others => '0');
    variable r257 : std_logic_vector(0 to 0) := (others => '0');
    variable r256 : std_logic_vector(0 to 0) := (others => '0');
    variable r255 : std_logic_vector(0 to 0) := (others => '0');
    variable r254 : std_logic_vector(0 to 0) := (others => '0');
    variable r253 : std_logic_vector(0 to 0) := (others => '0');
    variable r252 : std_logic_vector(0 to 0) := (others => '0');
    variable r251 : std_logic_vector(0 to 0) := (others => '0');
    variable r250 : std_logic_vector(0 to 0) := (others => '0');
    variable r249 : std_logic_vector(0 to 0) := (others => '0');
    variable r248 : std_logic_vector(0 to 0) := (others => '0');
    variable r247 : std_logic_vector(0 to 0) := (others => '0');
    variable r246 : std_logic_vector(0 to 0) := (others => '0');
    variable r245 : std_logic_vector(0 to 0) := (others => '0');
    variable r244 : std_logic_vector(0 to 0) := (others => '0');
    variable r243 : std_logic_vector(0 to 0) := (others => '0');
    variable r242 : std_logic_vector(0 to 0) := (others => '0');
    variable r241 : std_logic_vector(0 to 0) := (others => '0');
    variable r240 : std_logic_vector(0 to 0) := (others => '0');
    variable r239 : std_logic_vector(0 to 0) := (others => '0');
    variable r238 : std_logic_vector(0 to 0) := (others => '0');
    variable r237 : std_logic_vector(0 to 0) := (others => '0');
    variable r236 : std_logic_vector(0 to 0) := (others => '0');
    variable r235 : std_logic_vector(0 to 0) := (others => '0');
    variable r234 : std_logic_vector(0 to 0) := (others => '0');
    variable r233 : std_logic_vector(0 to 0) := (others => '0');
    variable r232 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r233 := "1";
    null;
    r234 := (r233);
    r235 := "0";
    null;
    r236 := (r235);
    r237 := "1";
    null;
    r238 := (r237);
    r239 := "0";
    null;
    r240 := (r239);
    r241 := "0";
    null;
    r242 := (r241);
    r243 := "1";
    null;
    r244 := (r243);
    r245 := "0";
    null;
    r246 := (r245);
    r247 := "1";
    null;
    r248 := (r247);
    r249 := "0";
    null;
    r250 := (r249);
    r251 := "1";
    null;
    r252 := (r251);
    r253 := "0";
    null;
    r254 := (r253);
    r255 := "0";
    null;
    r256 := (r255);
    r257 := "1";
    null;
    r258 := (r257);
    r259 := "1";
    null;
    r260 := (r259);
    r261 := "1";
    null;
    r262 := (r261);
    r263 := "1";
    null;
    r264 := (r263);
    r265 := "1";
    null;
    r266 := (r265);
    r267 := "1";
    null;
    r268 := (r267);
    r269 := "1";
    null;
    r270 := (r269);
    r271 := "1";
    null;
    r272 := (r271);
    r273 := "0";
    null;
    r274 := (r273);
    r275 := "1";
    null;
    r276 := (r275);
    r277 := "0";
    null;
    r278 := (r277);
    r279 := "1";
    null;
    r280 := (r279);
    r281 := "0";
    null;
    r282 := (r281);
    r283 := "0";
    null;
    r284 := (r283);
    r285 := "1";
    null;
    r286 := (r285);
    r287 := "1";
    null;
    r288 := (r287);
    r289 := "1";
    null;
    r290 := (r289);
    r291 := "0";
    null;
    r292 := (r291);
    r293 := "1";
    null;
    r294 := (r293);
    r295 := "0";
    null;
    r296 := (r295);
    r232 := (r234 & r236 & r238 & r240 & r242 & r244 & r246 & r248 & r250 & r252 & r254 & r256 & r258 & r260 & r262 & r264 & r266 & r268 & r270 & r272 & r274 & r276 & r278 & r280 & r282 & r284 & r286 & r288 & r290 & r292 & r294 & r296);
    return r232;
  end rewire_MetaprogrammingRWwa54ff53a_231;
  function rewire_MetaprogrammingRWw3c6ef372_164 return std_logic_vector
  is
    variable r229 : std_logic_vector(0 to 0) := (others => '0');
    variable r228 : std_logic_vector(0 to 0) := (others => '0');
    variable r227 : std_logic_vector(0 to 0) := (others => '0');
    variable r226 : std_logic_vector(0 to 0) := (others => '0');
    variable r225 : std_logic_vector(0 to 0) := (others => '0');
    variable r224 : std_logic_vector(0 to 0) := (others => '0');
    variable r223 : std_logic_vector(0 to 0) := (others => '0');
    variable r222 : std_logic_vector(0 to 0) := (others => '0');
    variable r221 : std_logic_vector(0 to 0) := (others => '0');
    variable r220 : std_logic_vector(0 to 0) := (others => '0');
    variable r219 : std_logic_vector(0 to 0) := (others => '0');
    variable r218 : std_logic_vector(0 to 0) := (others => '0');
    variable r217 : std_logic_vector(0 to 0) := (others => '0');
    variable r216 : std_logic_vector(0 to 0) := (others => '0');
    variable r215 : std_logic_vector(0 to 0) := (others => '0');
    variable r214 : std_logic_vector(0 to 0) := (others => '0');
    variable r213 : std_logic_vector(0 to 0) := (others => '0');
    variable r212 : std_logic_vector(0 to 0) := (others => '0');
    variable r211 : std_logic_vector(0 to 0) := (others => '0');
    variable r210 : std_logic_vector(0 to 0) := (others => '0');
    variable r209 : std_logic_vector(0 to 0) := (others => '0');
    variable r208 : std_logic_vector(0 to 0) := (others => '0');
    variable r207 : std_logic_vector(0 to 0) := (others => '0');
    variable r206 : std_logic_vector(0 to 0) := (others => '0');
    variable r205 : std_logic_vector(0 to 0) := (others => '0');
    variable r204 : std_logic_vector(0 to 0) := (others => '0');
    variable r203 : std_logic_vector(0 to 0) := (others => '0');
    variable r202 : std_logic_vector(0 to 0) := (others => '0');
    variable r201 : std_logic_vector(0 to 0) := (others => '0');
    variable r200 : std_logic_vector(0 to 0) := (others => '0');
    variable r199 : std_logic_vector(0 to 0) := (others => '0');
    variable r198 : std_logic_vector(0 to 0) := (others => '0');
    variable r197 : std_logic_vector(0 to 0) := (others => '0');
    variable r196 : std_logic_vector(0 to 0) := (others => '0');
    variable r195 : std_logic_vector(0 to 0) := (others => '0');
    variable r194 : std_logic_vector(0 to 0) := (others => '0');
    variable r193 : std_logic_vector(0 to 0) := (others => '0');
    variable r192 : std_logic_vector(0 to 0) := (others => '0');
    variable r191 : std_logic_vector(0 to 0) := (others => '0');
    variable r190 : std_logic_vector(0 to 0) := (others => '0');
    variable r189 : std_logic_vector(0 to 0) := (others => '0');
    variable r188 : std_logic_vector(0 to 0) := (others => '0');
    variable r187 : std_logic_vector(0 to 0) := (others => '0');
    variable r186 : std_logic_vector(0 to 0) := (others => '0');
    variable r185 : std_logic_vector(0 to 0) := (others => '0');
    variable r184 : std_logic_vector(0 to 0) := (others => '0');
    variable r183 : std_logic_vector(0 to 0) := (others => '0');
    variable r182 : std_logic_vector(0 to 0) := (others => '0');
    variable r181 : std_logic_vector(0 to 0) := (others => '0');
    variable r180 : std_logic_vector(0 to 0) := (others => '0');
    variable r179 : std_logic_vector(0 to 0) := (others => '0');
    variable r178 : std_logic_vector(0 to 0) := (others => '0');
    variable r177 : std_logic_vector(0 to 0) := (others => '0');
    variable r176 : std_logic_vector(0 to 0) := (others => '0');
    variable r175 : std_logic_vector(0 to 0) := (others => '0');
    variable r174 : std_logic_vector(0 to 0) := (others => '0');
    variable r173 : std_logic_vector(0 to 0) := (others => '0');
    variable r172 : std_logic_vector(0 to 0) := (others => '0');
    variable r171 : std_logic_vector(0 to 0) := (others => '0');
    variable r170 : std_logic_vector(0 to 0) := (others => '0');
    variable r169 : std_logic_vector(0 to 0) := (others => '0');
    variable r168 : std_logic_vector(0 to 0) := (others => '0');
    variable r167 : std_logic_vector(0 to 0) := (others => '0');
    variable r166 : std_logic_vector(0 to 0) := (others => '0');
    variable r165 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r166 := "0";
    null;
    r167 := (r166);
    r168 := "0";
    null;
    r169 := (r168);
    r170 := "1";
    null;
    r171 := (r170);
    r172 := "1";
    null;
    r173 := (r172);
    r174 := "1";
    null;
    r175 := (r174);
    r176 := "1";
    null;
    r177 := (r176);
    r178 := "0";
    null;
    r179 := (r178);
    r180 := "0";
    null;
    r181 := (r180);
    r182 := "0";
    null;
    r183 := (r182);
    r184 := "1";
    null;
    r185 := (r184);
    r186 := "1";
    null;
    r187 := (r186);
    r188 := "0";
    null;
    r189 := (r188);
    r190 := "1";
    null;
    r191 := (r190);
    r192 := "1";
    null;
    r193 := (r192);
    r194 := "1";
    null;
    r195 := (r194);
    r196 := "0";
    null;
    r197 := (r196);
    r198 := "1";
    null;
    r199 := (r198);
    r200 := "1";
    null;
    r201 := (r200);
    r202 := "1";
    null;
    r203 := (r202);
    r204 := "1";
    null;
    r205 := (r204);
    r206 := "0";
    null;
    r207 := (r206);
    r208 := "0";
    null;
    r209 := (r208);
    r210 := "1";
    null;
    r211 := (r210);
    r212 := "1";
    null;
    r213 := (r212);
    r214 := "0";
    null;
    r215 := (r214);
    r216 := "1";
    null;
    r217 := (r216);
    r218 := "1";
    null;
    r219 := (r218);
    r220 := "1";
    null;
    r221 := (r220);
    r222 := "0";
    null;
    r223 := (r222);
    r224 := "0";
    null;
    r225 := (r224);
    r226 := "1";
    null;
    r227 := (r226);
    r228 := "0";
    null;
    r229 := (r228);
    r165 := (r167 & r169 & r171 & r173 & r175 & r177 & r179 & r181 & r183 & r185 & r187 & r189 & r191 & r193 & r195 & r197 & r199 & r201 & r203 & r205 & r207 & r209 & r211 & r213 & r215 & r217 & r219 & r221 & r223 & r225 & r227 & r229);
    return r165;
  end rewire_MetaprogrammingRWw3c6ef372_164;
  function rewire_MetaprogrammingRWwbb67ae85_97 return std_logic_vector
  is
    variable r162 : std_logic_vector(0 to 0) := (others => '0');
    variable r161 : std_logic_vector(0 to 0) := (others => '0');
    variable r160 : std_logic_vector(0 to 0) := (others => '0');
    variable r159 : std_logic_vector(0 to 0) := (others => '0');
    variable r158 : std_logic_vector(0 to 0) := (others => '0');
    variable r157 : std_logic_vector(0 to 0) := (others => '0');
    variable r156 : std_logic_vector(0 to 0) := (others => '0');
    variable r155 : std_logic_vector(0 to 0) := (others => '0');
    variable r154 : std_logic_vector(0 to 0) := (others => '0');
    variable r153 : std_logic_vector(0 to 0) := (others => '0');
    variable r152 : std_logic_vector(0 to 0) := (others => '0');
    variable r151 : std_logic_vector(0 to 0) := (others => '0');
    variable r150 : std_logic_vector(0 to 0) := (others => '0');
    variable r149 : std_logic_vector(0 to 0) := (others => '0');
    variable r148 : std_logic_vector(0 to 0) := (others => '0');
    variable r147 : std_logic_vector(0 to 0) := (others => '0');
    variable r146 : std_logic_vector(0 to 0) := (others => '0');
    variable r145 : std_logic_vector(0 to 0) := (others => '0');
    variable r144 : std_logic_vector(0 to 0) := (others => '0');
    variable r143 : std_logic_vector(0 to 0) := (others => '0');
    variable r142 : std_logic_vector(0 to 0) := (others => '0');
    variable r141 : std_logic_vector(0 to 0) := (others => '0');
    variable r140 : std_logic_vector(0 to 0) := (others => '0');
    variable r139 : std_logic_vector(0 to 0) := (others => '0');
    variable r138 : std_logic_vector(0 to 0) := (others => '0');
    variable r137 : std_logic_vector(0 to 0) := (others => '0');
    variable r136 : std_logic_vector(0 to 0) := (others => '0');
    variable r135 : std_logic_vector(0 to 0) := (others => '0');
    variable r134 : std_logic_vector(0 to 0) := (others => '0');
    variable r133 : std_logic_vector(0 to 0) := (others => '0');
    variable r132 : std_logic_vector(0 to 0) := (others => '0');
    variable r131 : std_logic_vector(0 to 0) := (others => '0');
    variable r130 : std_logic_vector(0 to 0) := (others => '0');
    variable r129 : std_logic_vector(0 to 0) := (others => '0');
    variable r128 : std_logic_vector(0 to 0) := (others => '0');
    variable r127 : std_logic_vector(0 to 0) := (others => '0');
    variable r126 : std_logic_vector(0 to 0) := (others => '0');
    variable r125 : std_logic_vector(0 to 0) := (others => '0');
    variable r124 : std_logic_vector(0 to 0) := (others => '0');
    variable r123 : std_logic_vector(0 to 0) := (others => '0');
    variable r122 : std_logic_vector(0 to 0) := (others => '0');
    variable r121 : std_logic_vector(0 to 0) := (others => '0');
    variable r120 : std_logic_vector(0 to 0) := (others => '0');
    variable r119 : std_logic_vector(0 to 0) := (others => '0');
    variable r118 : std_logic_vector(0 to 0) := (others => '0');
    variable r117 : std_logic_vector(0 to 0) := (others => '0');
    variable r116 : std_logic_vector(0 to 0) := (others => '0');
    variable r115 : std_logic_vector(0 to 0) := (others => '0');
    variable r114 : std_logic_vector(0 to 0) := (others => '0');
    variable r113 : std_logic_vector(0 to 0) := (others => '0');
    variable r112 : std_logic_vector(0 to 0) := (others => '0');
    variable r111 : std_logic_vector(0 to 0) := (others => '0');
    variable r110 : std_logic_vector(0 to 0) := (others => '0');
    variable r109 : std_logic_vector(0 to 0) := (others => '0');
    variable r108 : std_logic_vector(0 to 0) := (others => '0');
    variable r107 : std_logic_vector(0 to 0) := (others => '0');
    variable r106 : std_logic_vector(0 to 0) := (others => '0');
    variable r105 : std_logic_vector(0 to 0) := (others => '0');
    variable r104 : std_logic_vector(0 to 0) := (others => '0');
    variable r103 : std_logic_vector(0 to 0) := (others => '0');
    variable r102 : std_logic_vector(0 to 0) := (others => '0');
    variable r101 : std_logic_vector(0 to 0) := (others => '0');
    variable r100 : std_logic_vector(0 to 0) := (others => '0');
    variable r99 : std_logic_vector(0 to 0) := (others => '0');
    variable r98 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r99 := "1";
    null;
    r100 := (r99);
    r101 := "0";
    null;
    r102 := (r101);
    r103 := "1";
    null;
    r104 := (r103);
    r105 := "1";
    null;
    r106 := (r105);
    r107 := "1";
    null;
    r108 := (r107);
    r109 := "0";
    null;
    r110 := (r109);
    r111 := "1";
    null;
    r112 := (r111);
    r113 := "1";
    null;
    r114 := (r113);
    r115 := "0";
    null;
    r116 := (r115);
    r117 := "1";
    null;
    r118 := (r117);
    r119 := "1";
    null;
    r120 := (r119);
    r121 := "0";
    null;
    r122 := (r121);
    r123 := "0";
    null;
    r124 := (r123);
    r125 := "1";
    null;
    r126 := (r125);
    r127 := "1";
    null;
    r128 := (r127);
    r129 := "1";
    null;
    r130 := (r129);
    r131 := "1";
    null;
    r132 := (r131);
    r133 := "0";
    null;
    r134 := (r133);
    r135 := "1";
    null;
    r136 := (r135);
    r137 := "0";
    null;
    r138 := (r137);
    r139 := "1";
    null;
    r140 := (r139);
    r141 := "1";
    null;
    r142 := (r141);
    r143 := "1";
    null;
    r144 := (r143);
    r145 := "0";
    null;
    r146 := (r145);
    r147 := "1";
    null;
    r148 := (r147);
    r149 := "0";
    null;
    r150 := (r149);
    r151 := "0";
    null;
    r152 := (r151);
    r153 := "0";
    null;
    r154 := (r153);
    r155 := "0";
    null;
    r156 := (r155);
    r157 := "1";
    null;
    r158 := (r157);
    r159 := "0";
    null;
    r160 := (r159);
    r161 := "1";
    null;
    r162 := (r161);
    r98 := (r100 & r102 & r104 & r106 & r108 & r110 & r112 & r114 & r116 & r118 & r120 & r122 & r124 & r126 & r128 & r130 & r132 & r134 & r136 & r138 & r140 & r142 & r144 & r146 & r148 & r150 & r152 & r154 & r156 & r158 & r160 & r162);
    return r98;
  end rewire_MetaprogrammingRWwbb67ae85_97;
  function rewire_MetaprogrammingRWw6a09e667_30 return std_logic_vector
  is
    variable r95 : std_logic_vector(0 to 0) := (others => '0');
    variable r94 : std_logic_vector(0 to 0) := (others => '0');
    variable r93 : std_logic_vector(0 to 0) := (others => '0');
    variable r92 : std_logic_vector(0 to 0) := (others => '0');
    variable r91 : std_logic_vector(0 to 0) := (others => '0');
    variable r90 : std_logic_vector(0 to 0) := (others => '0');
    variable r89 : std_logic_vector(0 to 0) := (others => '0');
    variable r88 : std_logic_vector(0 to 0) := (others => '0');
    variable r87 : std_logic_vector(0 to 0) := (others => '0');
    variable r86 : std_logic_vector(0 to 0) := (others => '0');
    variable r85 : std_logic_vector(0 to 0) := (others => '0');
    variable r84 : std_logic_vector(0 to 0) := (others => '0');
    variable r83 : std_logic_vector(0 to 0) := (others => '0');
    variable r82 : std_logic_vector(0 to 0) := (others => '0');
    variable r81 : std_logic_vector(0 to 0) := (others => '0');
    variable r80 : std_logic_vector(0 to 0) := (others => '0');
    variable r79 : std_logic_vector(0 to 0) := (others => '0');
    variable r78 : std_logic_vector(0 to 0) := (others => '0');
    variable r77 : std_logic_vector(0 to 0) := (others => '0');
    variable r76 : std_logic_vector(0 to 0) := (others => '0');
    variable r75 : std_logic_vector(0 to 0) := (others => '0');
    variable r74 : std_logic_vector(0 to 0) := (others => '0');
    variable r73 : std_logic_vector(0 to 0) := (others => '0');
    variable r72 : std_logic_vector(0 to 0) := (others => '0');
    variable r71 : std_logic_vector(0 to 0) := (others => '0');
    variable r70 : std_logic_vector(0 to 0) := (others => '0');
    variable r69 : std_logic_vector(0 to 0) := (others => '0');
    variable r68 : std_logic_vector(0 to 0) := (others => '0');
    variable r67 : std_logic_vector(0 to 0) := (others => '0');
    variable r66 : std_logic_vector(0 to 0) := (others => '0');
    variable r65 : std_logic_vector(0 to 0) := (others => '0');
    variable r64 : std_logic_vector(0 to 0) := (others => '0');
    variable r63 : std_logic_vector(0 to 0) := (others => '0');
    variable r62 : std_logic_vector(0 to 0) := (others => '0');
    variable r61 : std_logic_vector(0 to 0) := (others => '0');
    variable r60 : std_logic_vector(0 to 0) := (others => '0');
    variable r59 : std_logic_vector(0 to 0) := (others => '0');
    variable r58 : std_logic_vector(0 to 0) := (others => '0');
    variable r57 : std_logic_vector(0 to 0) := (others => '0');
    variable r56 : std_logic_vector(0 to 0) := (others => '0');
    variable r55 : std_logic_vector(0 to 0) := (others => '0');
    variable r54 : std_logic_vector(0 to 0) := (others => '0');
    variable r53 : std_logic_vector(0 to 0) := (others => '0');
    variable r52 : std_logic_vector(0 to 0) := (others => '0');
    variable r51 : std_logic_vector(0 to 0) := (others => '0');
    variable r50 : std_logic_vector(0 to 0) := (others => '0');
    variable r49 : std_logic_vector(0 to 0) := (others => '0');
    variable r48 : std_logic_vector(0 to 0) := (others => '0');
    variable r47 : std_logic_vector(0 to 0) := (others => '0');
    variable r46 : std_logic_vector(0 to 0) := (others => '0');
    variable r45 : std_logic_vector(0 to 0) := (others => '0');
    variable r44 : std_logic_vector(0 to 0) := (others => '0');
    variable r43 : std_logic_vector(0 to 0) := (others => '0');
    variable r42 : std_logic_vector(0 to 0) := (others => '0');
    variable r41 : std_logic_vector(0 to 0) := (others => '0');
    variable r40 : std_logic_vector(0 to 0) := (others => '0');
    variable r39 : std_logic_vector(0 to 0) := (others => '0');
    variable r38 : std_logic_vector(0 to 0) := (others => '0');
    variable r37 : std_logic_vector(0 to 0) := (others => '0');
    variable r36 : std_logic_vector(0 to 0) := (others => '0');
    variable r35 : std_logic_vector(0 to 0) := (others => '0');
    variable r34 : std_logic_vector(0 to 0) := (others => '0');
    variable r33 : std_logic_vector(0 to 0) := (others => '0');
    variable r32 : std_logic_vector(0 to 0) := (others => '0');
    variable r31 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r32 := "0";
    null;
    r33 := (r32);
    r34 := "1";
    null;
    r35 := (r34);
    r36 := "1";
    null;
    r37 := (r36);
    r38 := "0";
    null;
    r39 := (r38);
    r40 := "1";
    null;
    r41 := (r40);
    r42 := "0";
    null;
    r43 := (r42);
    r44 := "1";
    null;
    r45 := (r44);
    r46 := "0";
    null;
    r47 := (r46);
    r48 := "0";
    null;
    r49 := (r48);
    r50 := "0";
    null;
    r51 := (r50);
    r52 := "0";
    null;
    r53 := (r52);
    r54 := "0";
    null;
    r55 := (r54);
    r56 := "1";
    null;
    r57 := (r56);
    r58 := "0";
    null;
    r59 := (r58);
    r60 := "0";
    null;
    r61 := (r60);
    r62 := "1";
    null;
    r63 := (r62);
    r64 := "1";
    null;
    r65 := (r64);
    r66 := "1";
    null;
    r67 := (r66);
    r68 := "1";
    null;
    r69 := (r68);
    r70 := "0";
    null;
    r71 := (r70);
    r72 := "0";
    null;
    r73 := (r72);
    r74 := "1";
    null;
    r75 := (r74);
    r76 := "1";
    null;
    r77 := (r76);
    r78 := "0";
    null;
    r79 := (r78);
    r80 := "0";
    null;
    r81 := (r80);
    r82 := "1";
    null;
    r83 := (r82);
    r84 := "1";
    null;
    r85 := (r84);
    r86 := "0";
    null;
    r87 := (r86);
    r88 := "0";
    null;
    r89 := (r88);
    r90 := "1";
    null;
    r91 := (r90);
    r92 := "1";
    null;
    r93 := (r92);
    r94 := "1";
    null;
    r95 := (r94);
    r31 := (r33 & r35 & r37 & r39 & r41 & r43 & r45 & r47 & r49 & r51 & r53 & r55 & r57 & r59 & r61 & r63 & r65 & r67 & r69 & r71 & r73 & r75 & r77 & r79 & r81 & r83 & r85 & r87 & r89 & r91 & r93 & r95);
    return r31;
  end rewire_MetaprogrammingRWw6a09e667_30;
  signal control_flop : control_state := STATE0;
  signal control_flop_next : control_state := STATE0;
  signal input_flop : std_logic_vector(0 to 67) := (others => '0');
  signal goto_L7851_flop : boolean := false;
  signal goto_L7844_flop : boolean := false;
  signal goto_L7806_flop : boolean := false;
  signal goto_L7767_flop : boolean := false;
  signal goto_L7728_flop : boolean := false;
  signal goto_L7570_flop : boolean := false;
  signal goto_L7690_flop : boolean := false;
  signal goto_L7575_flop : boolean := false;
  signal goto_L1784_flop : boolean := false;
  signal goto_L1785_flop : boolean := false;
  signal goto_L1638_flop : boolean := false;
  signal goto_L1502_flop : boolean := false;
  signal goto_L1366_flop : boolean := false;
  signal goto_L1230_flop : boolean := false;
  signal goto_L1094_flop : boolean := false;
  signal goto_L958_flop : boolean := false;
  signal goto_L822_flop : boolean := false;
  signal goto_L686_flop : boolean := false;
  signal goto_L11_flop : boolean := false;
  signal goto_L13_flop : boolean := false;
  signal goto_L690_flop : boolean := false;
  signal goto_L826_flop : boolean := false;
  signal goto_L962_flop : boolean := false;
  signal goto_L1098_flop : boolean := false;
  signal goto_L1234_flop : boolean := false;
  signal goto_L1370_flop : boolean := false;
  signal goto_L1506_flop : boolean := false;
  signal goto_L1642_flop : boolean := false;
  signal goto_L7693_flop : boolean := false;
  signal goto_L7732_flop : boolean := false;
  signal goto_L7771_flop : boolean := false;
  signal goto_L7810_flop : boolean := false;
  signal goto_L7777_flop : boolean := false;
  signal goto_L7738_flop : boolean := false;
  signal goto_L7699_flop : boolean := false;
  signal goto_L1658_flop : boolean := false;
  signal goto_L1522_flop : boolean := false;
  signal goto_L1386_flop : boolean := false;
  signal goto_L1250_flop : boolean := false;
  signal goto_L1114_flop : boolean := false;
  signal goto_L978_flop : boolean := false;
  signal goto_L842_flop : boolean := false;
  signal goto_L706_flop : boolean := false;
  signal goto_L567_flop : boolean := false;
  signal goto_L0_flop : boolean := false;
  signal goto_L7852_flop : boolean := false;
  signal r7843_flop : std_logic_vector(0 to 67) := (others => '0');
  signal r7840_flop : std_logic_vector(0 to 64) := (others => '0');
  signal r7817_flop : std_logic_vector(0 to 255) := (others => '0');
  signal r7814_flop : std_logic_vector(0 to 255) := (others => '0');
  signal r7805_flop : std_logic_vector(0 to 67) := (others => '0');
  signal r7802_flop : std_logic_vector(0 to 64) := (others => '0');
  signal r7779_flop : std_logic_vector(0 to 255) := (others => '0');
  signal r7776_flop : std_logic_vector(0 to 255) := (others => '0');
  signal b7774_flop : boolean := false;
  signal r7766_flop : std_logic_vector(0 to 67) := (others => '0');
  signal r7763_flop : std_logic_vector(0 to 64) := (others => '0');
  signal r7740_flop : std_logic_vector(0 to 255) := (others => '0');
  signal r7737_flop : std_logic_vector(0 to 255) := (others => '0');
  signal b7735_flop : boolean := false;
  signal r7727_flop : std_logic_vector(0 to 67) := (others => '0');
  signal r7724_flop : std_logic_vector(0 to 64) := (others => '0');
  signal r7701_flop : std_logic_vector(0 to 255) := (others => '0');
  signal r7698_flop : std_logic_vector(0 to 255) := (others => '0');
  signal b7696_flop : boolean := false;
  signal r7679_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r7675_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r7671_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r7667_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r7663_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r7659_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r7655_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r7651_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r7647_flop : std_logic_vector(0 to 255) := (others => '0');
  signal b7644_flop : boolean := false;
  signal b7642_flop : boolean := false;
  signal b7640_flop : boolean := false;
  signal b7638_flop : boolean := false;
  signal b7636_flop : boolean := false;
  signal b7634_flop : boolean := false;
  signal b7632_flop : boolean := false;
  signal b7630_flop : boolean := false;
  signal r7628_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r7626_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r7624_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r7622_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r7620_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r7618_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r7616_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r7614_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r7610_flop : std_logic_vector(0 to 255) := (others => '0');
  signal b7608_flop : boolean := false;
  signal b7606_flop : boolean := false;
  signal b7604_flop : boolean := false;
  signal b7602_flop : boolean := false;
  signal b7600_flop : boolean := false;
  signal b7598_flop : boolean := false;
  signal b7596_flop : boolean := false;
  signal b7594_flop : boolean := false;
  signal r7592_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r7590_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r7588_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r7586_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r7584_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r7582_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r7580_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r7578_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r7574_flop : std_logic_vector(0 to 255) := (others => '0');
  signal b7572_flop : boolean := false;
  signal r7569_flop : std_logic_vector(0 to 67) := (others => '0');
  signal r7565_flop : std_logic_vector(0 to 63) := (others => '0');
  signal r7564_flop : std_logic_vector(0 to 64) := (others => '0');
  signal r7562_flop : std_logic_vector(0 to 0) := (others => '0');
  signal r7558_flop : std_logic_vector(0 to 5) := (others => '0');
  signal r7300_flop : std_logic_vector(0 to 5) := (others => '0');
  signal r7296_flop : std_logic_vector(0 to 255) := (others => '0');
  signal r7292_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r2874_flop : std_logic_vector(0 to 5) := (others => '0');
  signal r2376_flop : std_logic_vector(0 to 255) := (others => '0');
  signal r2375_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r2374_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r2371_flop : std_logic_vector(0 to 255) := (others => '0');
  signal r2365_flop : std_logic_vector(0 to 511) := (others => '0');
  signal r1862_flop : std_logic_vector(0 to 511) := (others => '0');
  signal b1859_flop : boolean := false;
  signal b1857_flop : boolean := false;
  signal b1855_flop : boolean := false;
  signal b1853_flop : boolean := false;
  signal b1851_flop : boolean := false;
  signal b1849_flop : boolean := false;
  signal b1847_flop : boolean := false;
  signal b1845_flop : boolean := false;
  signal b1843_flop : boolean := false;
  signal b1841_flop : boolean := false;
  signal b1839_flop : boolean := false;
  signal b1837_flop : boolean := false;
  signal b1835_flop : boolean := false;
  signal b1833_flop : boolean := false;
  signal b1831_flop : boolean := false;
  signal b1829_flop : boolean := false;
  signal r1827_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1825_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1823_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1821_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1819_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1817_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1815_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1813_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1811_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1809_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1807_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1805_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1803_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1801_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1799_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1797_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1795_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1792_flop : std_logic_vector(0 to 511) := (others => '0');
  signal r1790_flop : std_logic_vector(0 to 5) := (others => '0');
  signal r1787_flop : std_logic_vector(0 to 5) := (others => '0');
  signal r1783_flop : std_logic_vector(0 to 67) := (others => '0');
  signal r1779_flop : std_logic_vector(0 to 63) := (others => '0');
  signal r1778_flop : std_logic_vector(0 to 64) := (others => '0');
  signal r1776_flop : std_logic_vector(0 to 0) := (others => '0');
  signal r1754_flop : std_logic_vector(0 to 511) := (others => '0');
  signal b1751_flop : boolean := false;
  signal b1749_flop : boolean := false;
  signal b1747_flop : boolean := false;
  signal b1745_flop : boolean := false;
  signal b1743_flop : boolean := false;
  signal b1741_flop : boolean := false;
  signal b1739_flop : boolean := false;
  signal b1737_flop : boolean := false;
  signal b1735_flop : boolean := false;
  signal b1733_flop : boolean := false;
  signal b1731_flop : boolean := false;
  signal b1729_flop : boolean := false;
  signal b1727_flop : boolean := false;
  signal b1725_flop : boolean := false;
  signal b1723_flop : boolean := false;
  signal b1721_flop : boolean := false;
  signal r1719_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1717_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1715_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1713_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1711_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1709_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1707_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1705_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1703_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1701_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1699_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1697_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1695_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1693_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1691_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1689_flop : std_logic_vector(0 to 31) := (others => '0');
  signal b1686_flop : boolean := false;
  signal b1684_flop : boolean := false;
  signal r1682_flop : std_logic_vector(0 to 511) := (others => '0');
  signal r1680_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1678_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1676_flop : std_logic_vector(0 to 511) := (others => '0');
  signal r1670_flop : std_logic_vector(0 to 575) := (others => '0');
  signal r1667_flop : std_logic_vector(0 to 511) := (others => '0');
  signal r1663_flop : std_logic_vector(0 to 255) := (others => '0');
  signal r1659_flop : std_logic_vector(0 to 5) := (others => '0');
  signal r1657_flop : std_logic_vector(0 to 5) := (others => '0');
  signal b1655_flop : boolean := false;
  signal b1653_flop : boolean := false;
  signal b1651_flop : boolean := false;
  signal r1649_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1647_flop : std_logic_vector(0 to 31) := (others => '0');
  signal b1645_flop : boolean := false;
  signal r1637_flop : std_logic_vector(0 to 67) := (others => '0');
  signal r1633_flop : std_logic_vector(0 to 63) := (others => '0');
  signal r1632_flop : std_logic_vector(0 to 64) := (others => '0');
  signal r1630_flop : std_logic_vector(0 to 0) := (others => '0');
  signal r1608_flop : std_logic_vector(0 to 511) := (others => '0');
  signal b1605_flop : boolean := false;
  signal b1603_flop : boolean := false;
  signal b1601_flop : boolean := false;
  signal b1599_flop : boolean := false;
  signal b1597_flop : boolean := false;
  signal b1595_flop : boolean := false;
  signal b1593_flop : boolean := false;
  signal b1591_flop : boolean := false;
  signal b1589_flop : boolean := false;
  signal b1587_flop : boolean := false;
  signal b1585_flop : boolean := false;
  signal b1583_flop : boolean := false;
  signal b1581_flop : boolean := false;
  signal b1579_flop : boolean := false;
  signal b1577_flop : boolean := false;
  signal b1575_flop : boolean := false;
  signal r1573_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1571_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1569_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1567_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1565_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1563_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1561_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1559_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1557_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1555_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1553_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1551_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1549_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1547_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1545_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1543_flop : std_logic_vector(0 to 31) := (others => '0');
  signal b1540_flop : boolean := false;
  signal b1538_flop : boolean := false;
  signal r1536_flop : std_logic_vector(0 to 511) := (others => '0');
  signal r1534_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1532_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1530_flop : std_logic_vector(0 to 511) := (others => '0');
  signal r1524_flop : std_logic_vector(0 to 575) := (others => '0');
  signal r1521_flop : std_logic_vector(0 to 511) := (others => '0');
  signal b1519_flop : boolean := false;
  signal b1517_flop : boolean := false;
  signal b1515_flop : boolean := false;
  signal r1513_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1511_flop : std_logic_vector(0 to 31) := (others => '0');
  signal b1509_flop : boolean := false;
  signal r1501_flop : std_logic_vector(0 to 67) := (others => '0');
  signal r1497_flop : std_logic_vector(0 to 63) := (others => '0');
  signal r1496_flop : std_logic_vector(0 to 64) := (others => '0');
  signal r1494_flop : std_logic_vector(0 to 0) := (others => '0');
  signal r1472_flop : std_logic_vector(0 to 511) := (others => '0');
  signal b1469_flop : boolean := false;
  signal b1467_flop : boolean := false;
  signal b1465_flop : boolean := false;
  signal b1463_flop : boolean := false;
  signal b1461_flop : boolean := false;
  signal b1459_flop : boolean := false;
  signal b1457_flop : boolean := false;
  signal b1455_flop : boolean := false;
  signal b1453_flop : boolean := false;
  signal b1451_flop : boolean := false;
  signal b1449_flop : boolean := false;
  signal b1447_flop : boolean := false;
  signal b1445_flop : boolean := false;
  signal b1443_flop : boolean := false;
  signal b1441_flop : boolean := false;
  signal b1439_flop : boolean := false;
  signal r1437_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1435_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1433_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1431_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1429_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1427_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1425_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1423_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1421_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1419_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1417_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1415_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1413_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1411_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1409_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1407_flop : std_logic_vector(0 to 31) := (others => '0');
  signal b1404_flop : boolean := false;
  signal b1402_flop : boolean := false;
  signal r1400_flop : std_logic_vector(0 to 511) := (others => '0');
  signal r1398_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1396_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1394_flop : std_logic_vector(0 to 511) := (others => '0');
  signal r1388_flop : std_logic_vector(0 to 575) := (others => '0');
  signal r1385_flop : std_logic_vector(0 to 511) := (others => '0');
  signal b1383_flop : boolean := false;
  signal b1381_flop : boolean := false;
  signal b1379_flop : boolean := false;
  signal r1377_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1375_flop : std_logic_vector(0 to 31) := (others => '0');
  signal b1373_flop : boolean := false;
  signal r1365_flop : std_logic_vector(0 to 67) := (others => '0');
  signal r1361_flop : std_logic_vector(0 to 63) := (others => '0');
  signal r1360_flop : std_logic_vector(0 to 64) := (others => '0');
  signal r1358_flop : std_logic_vector(0 to 0) := (others => '0');
  signal r1336_flop : std_logic_vector(0 to 511) := (others => '0');
  signal b1333_flop : boolean := false;
  signal b1331_flop : boolean := false;
  signal b1329_flop : boolean := false;
  signal b1327_flop : boolean := false;
  signal b1325_flop : boolean := false;
  signal b1323_flop : boolean := false;
  signal b1321_flop : boolean := false;
  signal b1319_flop : boolean := false;
  signal b1317_flop : boolean := false;
  signal b1315_flop : boolean := false;
  signal b1313_flop : boolean := false;
  signal b1311_flop : boolean := false;
  signal b1309_flop : boolean := false;
  signal b1307_flop : boolean := false;
  signal b1305_flop : boolean := false;
  signal b1303_flop : boolean := false;
  signal r1301_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1299_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1297_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1295_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1293_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1291_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1289_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1287_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1285_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1283_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1281_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1279_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1277_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1275_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1273_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1271_flop : std_logic_vector(0 to 31) := (others => '0');
  signal b1268_flop : boolean := false;
  signal b1266_flop : boolean := false;
  signal r1264_flop : std_logic_vector(0 to 511) := (others => '0');
  signal r1262_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1260_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1258_flop : std_logic_vector(0 to 511) := (others => '0');
  signal r1252_flop : std_logic_vector(0 to 575) := (others => '0');
  signal r1249_flop : std_logic_vector(0 to 511) := (others => '0');
  signal b1247_flop : boolean := false;
  signal b1245_flop : boolean := false;
  signal b1243_flop : boolean := false;
  signal r1241_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1239_flop : std_logic_vector(0 to 31) := (others => '0');
  signal b1237_flop : boolean := false;
  signal r1229_flop : std_logic_vector(0 to 67) := (others => '0');
  signal r1225_flop : std_logic_vector(0 to 63) := (others => '0');
  signal r1224_flop : std_logic_vector(0 to 64) := (others => '0');
  signal r1222_flop : std_logic_vector(0 to 0) := (others => '0');
  signal r1200_flop : std_logic_vector(0 to 511) := (others => '0');
  signal b1197_flop : boolean := false;
  signal b1195_flop : boolean := false;
  signal b1193_flop : boolean := false;
  signal b1191_flop : boolean := false;
  signal b1189_flop : boolean := false;
  signal b1187_flop : boolean := false;
  signal b1185_flop : boolean := false;
  signal b1183_flop : boolean := false;
  signal b1181_flop : boolean := false;
  signal b1179_flop : boolean := false;
  signal b1177_flop : boolean := false;
  signal b1175_flop : boolean := false;
  signal b1173_flop : boolean := false;
  signal b1171_flop : boolean := false;
  signal b1169_flop : boolean := false;
  signal b1167_flop : boolean := false;
  signal r1165_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1163_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1161_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1159_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1157_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1155_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1153_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1151_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1149_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1147_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1145_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1143_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1141_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1139_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1137_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1135_flop : std_logic_vector(0 to 31) := (others => '0');
  signal b1132_flop : boolean := false;
  signal b1130_flop : boolean := false;
  signal r1128_flop : std_logic_vector(0 to 511) := (others => '0');
  signal r1126_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1124_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1122_flop : std_logic_vector(0 to 511) := (others => '0');
  signal r1116_flop : std_logic_vector(0 to 575) := (others => '0');
  signal r1113_flop : std_logic_vector(0 to 511) := (others => '0');
  signal b1111_flop : boolean := false;
  signal b1109_flop : boolean := false;
  signal b1107_flop : boolean := false;
  signal r1105_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1103_flop : std_logic_vector(0 to 31) := (others => '0');
  signal b1101_flop : boolean := false;
  signal r1093_flop : std_logic_vector(0 to 67) := (others => '0');
  signal r1089_flop : std_logic_vector(0 to 63) := (others => '0');
  signal r1088_flop : std_logic_vector(0 to 64) := (others => '0');
  signal r1086_flop : std_logic_vector(0 to 0) := (others => '0');
  signal r1064_flop : std_logic_vector(0 to 511) := (others => '0');
  signal b1061_flop : boolean := false;
  signal b1059_flop : boolean := false;
  signal b1057_flop : boolean := false;
  signal b1055_flop : boolean := false;
  signal b1053_flop : boolean := false;
  signal b1051_flop : boolean := false;
  signal b1049_flop : boolean := false;
  signal b1047_flop : boolean := false;
  signal b1045_flop : boolean := false;
  signal b1043_flop : boolean := false;
  signal b1041_flop : boolean := false;
  signal b1039_flop : boolean := false;
  signal b1037_flop : boolean := false;
  signal b1035_flop : boolean := false;
  signal b1033_flop : boolean := false;
  signal b1031_flop : boolean := false;
  signal r1029_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1027_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1025_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1023_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1021_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1019_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1017_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1015_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1013_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1011_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1009_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1007_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1005_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1003_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1001_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r999_flop : std_logic_vector(0 to 31) := (others => '0');
  signal b996_flop : boolean := false;
  signal b994_flop : boolean := false;
  signal r992_flop : std_logic_vector(0 to 511) := (others => '0');
  signal r990_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r988_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r986_flop : std_logic_vector(0 to 511) := (others => '0');
  signal r980_flop : std_logic_vector(0 to 575) := (others => '0');
  signal r977_flop : std_logic_vector(0 to 511) := (others => '0');
  signal b975_flop : boolean := false;
  signal b973_flop : boolean := false;
  signal b971_flop : boolean := false;
  signal r969_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r967_flop : std_logic_vector(0 to 31) := (others => '0');
  signal b965_flop : boolean := false;
  signal r957_flop : std_logic_vector(0 to 67) := (others => '0');
  signal r953_flop : std_logic_vector(0 to 63) := (others => '0');
  signal r952_flop : std_logic_vector(0 to 64) := (others => '0');
  signal r950_flop : std_logic_vector(0 to 0) := (others => '0');
  signal r928_flop : std_logic_vector(0 to 511) := (others => '0');
  signal b925_flop : boolean := false;
  signal b923_flop : boolean := false;
  signal b921_flop : boolean := false;
  signal b919_flop : boolean := false;
  signal b917_flop : boolean := false;
  signal b915_flop : boolean := false;
  signal b913_flop : boolean := false;
  signal b911_flop : boolean := false;
  signal b909_flop : boolean := false;
  signal b907_flop : boolean := false;
  signal b905_flop : boolean := false;
  signal b903_flop : boolean := false;
  signal b901_flop : boolean := false;
  signal b899_flop : boolean := false;
  signal b897_flop : boolean := false;
  signal b895_flop : boolean := false;
  signal r893_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r891_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r889_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r887_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r885_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r883_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r881_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r879_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r877_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r875_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r873_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r871_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r869_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r867_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r865_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r863_flop : std_logic_vector(0 to 31) := (others => '0');
  signal b860_flop : boolean := false;
  signal b858_flop : boolean := false;
  signal r856_flop : std_logic_vector(0 to 511) := (others => '0');
  signal r854_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r852_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r850_flop : std_logic_vector(0 to 511) := (others => '0');
  signal r844_flop : std_logic_vector(0 to 575) := (others => '0');
  signal r841_flop : std_logic_vector(0 to 511) := (others => '0');
  signal b839_flop : boolean := false;
  signal b837_flop : boolean := false;
  signal b835_flop : boolean := false;
  signal r833_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r831_flop : std_logic_vector(0 to 31) := (others => '0');
  signal b829_flop : boolean := false;
  signal r821_flop : std_logic_vector(0 to 67) := (others => '0');
  signal r817_flop : std_logic_vector(0 to 63) := (others => '0');
  signal r816_flop : std_logic_vector(0 to 64) := (others => '0');
  signal r814_flop : std_logic_vector(0 to 0) := (others => '0');
  signal r792_flop : std_logic_vector(0 to 511) := (others => '0');
  signal b789_flop : boolean := false;
  signal b787_flop : boolean := false;
  signal b785_flop : boolean := false;
  signal b783_flop : boolean := false;
  signal b781_flop : boolean := false;
  signal b779_flop : boolean := false;
  signal b777_flop : boolean := false;
  signal b775_flop : boolean := false;
  signal b773_flop : boolean := false;
  signal b771_flop : boolean := false;
  signal b769_flop : boolean := false;
  signal b767_flop : boolean := false;
  signal b765_flop : boolean := false;
  signal b763_flop : boolean := false;
  signal b761_flop : boolean := false;
  signal b759_flop : boolean := false;
  signal r757_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r755_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r753_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r751_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r749_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r747_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r745_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r743_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r741_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r739_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r737_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r735_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r733_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r731_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r729_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r727_flop : std_logic_vector(0 to 31) := (others => '0');
  signal b724_flop : boolean := false;
  signal b722_flop : boolean := false;
  signal r720_flop : std_logic_vector(0 to 511) := (others => '0');
  signal r718_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r716_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r714_flop : std_logic_vector(0 to 511) := (others => '0');
  signal r708_flop : std_logic_vector(0 to 575) := (others => '0');
  signal r705_flop : std_logic_vector(0 to 511) := (others => '0');
  signal b703_flop : boolean := false;
  signal b701_flop : boolean := false;
  signal b699_flop : boolean := false;
  signal r697_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r695_flop : std_logic_vector(0 to 31) := (others => '0');
  signal b693_flop : boolean := false;
  signal r685_flop : std_logic_vector(0 to 67) := (others => '0');
  signal r681_flop : std_logic_vector(0 to 63) := (others => '0');
  signal r680_flop : std_logic_vector(0 to 64) := (others => '0');
  signal r678_flop : std_logic_vector(0 to 0) := (others => '0');
  signal r656_flop : std_logic_vector(0 to 511) := (others => '0');
  signal b653_flop : boolean := false;
  signal b651_flop : boolean := false;
  signal b649_flop : boolean := false;
  signal b647_flop : boolean := false;
  signal b645_flop : boolean := false;
  signal b643_flop : boolean := false;
  signal b641_flop : boolean := false;
  signal b639_flop : boolean := false;
  signal b637_flop : boolean := false;
  signal b635_flop : boolean := false;
  signal b633_flop : boolean := false;
  signal b631_flop : boolean := false;
  signal b629_flop : boolean := false;
  signal b627_flop : boolean := false;
  signal b625_flop : boolean := false;
  signal b623_flop : boolean := false;
  signal r621_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r619_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r617_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r615_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r613_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r611_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r609_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r607_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r605_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r603_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r601_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r599_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r597_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r595_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r593_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r591_flop : std_logic_vector(0 to 31) := (others => '0');
  signal b588_flop : boolean := false;
  signal b586_flop : boolean := false;
  signal r584_flop : std_logic_vector(0 to 511) := (others => '0');
  signal r582_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r580_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r578_flop : std_logic_vector(0 to 511) := (others => '0');
  signal r572_flop : std_logic_vector(0 to 575) := (others => '0');
  signal r569_flop : std_logic_vector(0 to 511) := (others => '0');
  signal r566_flop : std_logic_vector(0 to 255) := (others => '0');
  signal b26_flop : boolean := false;
  signal b24_flop : boolean := false;
  signal b22_flop : boolean := false;
  signal r20_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r18_flop : std_logic_vector(0 to 31) := (others => '0');
  signal b16_flop : boolean := false;
  signal r12_flop : std_logic_vector(0 to 67) := (others => '0');
  signal r10_flop : std_logic_vector(0 to 67) := (others => '0');
  signal r6_flop : std_logic_vector(0 to 63) := (others => '0');
  signal r5_flop : std_logic_vector(0 to 64) := (others => '0');
  signal r3_flop : std_logic_vector(0 to 0) := (others => '0');
  signal statevar0_flop : std_logic_vector(0 to 255) := (others => '0');
  signal statevar1_flop : std_logic_vector(0 to 511) := (others => '0');
  signal statevar2_flop : std_logic_vector(0 to 255) := (others => '0');
  signal statevar3_flop : std_logic_vector(0 to 5) := (others => '0');
  signal goto_L7851_flop_next : boolean := false;
  signal goto_L7844_flop_next : boolean := false;
  signal goto_L7806_flop_next : boolean := false;
  signal goto_L7767_flop_next : boolean := false;
  signal goto_L7728_flop_next : boolean := false;
  signal goto_L7570_flop_next : boolean := false;
  signal goto_L7690_flop_next : boolean := false;
  signal goto_L7575_flop_next : boolean := false;
  signal goto_L1784_flop_next : boolean := false;
  signal goto_L1785_flop_next : boolean := false;
  signal goto_L1638_flop_next : boolean := false;
  signal goto_L1502_flop_next : boolean := false;
  signal goto_L1366_flop_next : boolean := false;
  signal goto_L1230_flop_next : boolean := false;
  signal goto_L1094_flop_next : boolean := false;
  signal goto_L958_flop_next : boolean := false;
  signal goto_L822_flop_next : boolean := false;
  signal goto_L686_flop_next : boolean := false;
  signal goto_L11_flop_next : boolean := false;
  signal goto_L13_flop_next : boolean := false;
  signal goto_L690_flop_next : boolean := false;
  signal goto_L826_flop_next : boolean := false;
  signal goto_L962_flop_next : boolean := false;
  signal goto_L1098_flop_next : boolean := false;
  signal goto_L1234_flop_next : boolean := false;
  signal goto_L1370_flop_next : boolean := false;
  signal goto_L1506_flop_next : boolean := false;
  signal goto_L1642_flop_next : boolean := false;
  signal goto_L7693_flop_next : boolean := false;
  signal goto_L7732_flop_next : boolean := false;
  signal goto_L7771_flop_next : boolean := false;
  signal goto_L7810_flop_next : boolean := false;
  signal goto_L7777_flop_next : boolean := false;
  signal goto_L7738_flop_next : boolean := false;
  signal goto_L7699_flop_next : boolean := false;
  signal goto_L1658_flop_next : boolean := false;
  signal goto_L1522_flop_next : boolean := false;
  signal goto_L1386_flop_next : boolean := false;
  signal goto_L1250_flop_next : boolean := false;
  signal goto_L1114_flop_next : boolean := false;
  signal goto_L978_flop_next : boolean := false;
  signal goto_L842_flop_next : boolean := false;
  signal goto_L706_flop_next : boolean := false;
  signal goto_L567_flop_next : boolean := false;
  signal goto_L0_flop_next : boolean := false;
  signal goto_L7852_flop_next : boolean := false;
  signal r7843_flop_next : std_logic_vector(0 to 67) := (others => '0');
  signal r7840_flop_next : std_logic_vector(0 to 64) := (others => '0');
  signal r7817_flop_next : std_logic_vector(0 to 255) := (others => '0');
  signal r7814_flop_next : std_logic_vector(0 to 255) := (others => '0');
  signal r7805_flop_next : std_logic_vector(0 to 67) := (others => '0');
  signal r7802_flop_next : std_logic_vector(0 to 64) := (others => '0');
  signal r7779_flop_next : std_logic_vector(0 to 255) := (others => '0');
  signal r7776_flop_next : std_logic_vector(0 to 255) := (others => '0');
  signal b7774_flop_next : boolean := false;
  signal r7766_flop_next : std_logic_vector(0 to 67) := (others => '0');
  signal r7763_flop_next : std_logic_vector(0 to 64) := (others => '0');
  signal r7740_flop_next : std_logic_vector(0 to 255) := (others => '0');
  signal r7737_flop_next : std_logic_vector(0 to 255) := (others => '0');
  signal b7735_flop_next : boolean := false;
  signal r7727_flop_next : std_logic_vector(0 to 67) := (others => '0');
  signal r7724_flop_next : std_logic_vector(0 to 64) := (others => '0');
  signal r7701_flop_next : std_logic_vector(0 to 255) := (others => '0');
  signal r7698_flop_next : std_logic_vector(0 to 255) := (others => '0');
  signal b7696_flop_next : boolean := false;
  signal r7679_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r7675_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r7671_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r7667_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r7663_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r7659_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r7655_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r7651_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r7647_flop_next : std_logic_vector(0 to 255) := (others => '0');
  signal b7644_flop_next : boolean := false;
  signal b7642_flop_next : boolean := false;
  signal b7640_flop_next : boolean := false;
  signal b7638_flop_next : boolean := false;
  signal b7636_flop_next : boolean := false;
  signal b7634_flop_next : boolean := false;
  signal b7632_flop_next : boolean := false;
  signal b7630_flop_next : boolean := false;
  signal r7628_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r7626_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r7624_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r7622_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r7620_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r7618_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r7616_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r7614_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r7610_flop_next : std_logic_vector(0 to 255) := (others => '0');
  signal b7608_flop_next : boolean := false;
  signal b7606_flop_next : boolean := false;
  signal b7604_flop_next : boolean := false;
  signal b7602_flop_next : boolean := false;
  signal b7600_flop_next : boolean := false;
  signal b7598_flop_next : boolean := false;
  signal b7596_flop_next : boolean := false;
  signal b7594_flop_next : boolean := false;
  signal r7592_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r7590_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r7588_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r7586_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r7584_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r7582_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r7580_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r7578_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r7574_flop_next : std_logic_vector(0 to 255) := (others => '0');
  signal b7572_flop_next : boolean := false;
  signal r7569_flop_next : std_logic_vector(0 to 67) := (others => '0');
  signal r7565_flop_next : std_logic_vector(0 to 63) := (others => '0');
  signal r7564_flop_next : std_logic_vector(0 to 64) := (others => '0');
  signal r7562_flop_next : std_logic_vector(0 to 0) := (others => '0');
  signal r7558_flop_next : std_logic_vector(0 to 5) := (others => '0');
  signal r7300_flop_next : std_logic_vector(0 to 5) := (others => '0');
  signal r7296_flop_next : std_logic_vector(0 to 255) := (others => '0');
  signal r7292_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r2874_flop_next : std_logic_vector(0 to 5) := (others => '0');
  signal r2376_flop_next : std_logic_vector(0 to 255) := (others => '0');
  signal r2375_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r2374_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r2371_flop_next : std_logic_vector(0 to 255) := (others => '0');
  signal r2365_flop_next : std_logic_vector(0 to 511) := (others => '0');
  signal r1862_flop_next : std_logic_vector(0 to 511) := (others => '0');
  signal b1859_flop_next : boolean := false;
  signal b1857_flop_next : boolean := false;
  signal b1855_flop_next : boolean := false;
  signal b1853_flop_next : boolean := false;
  signal b1851_flop_next : boolean := false;
  signal b1849_flop_next : boolean := false;
  signal b1847_flop_next : boolean := false;
  signal b1845_flop_next : boolean := false;
  signal b1843_flop_next : boolean := false;
  signal b1841_flop_next : boolean := false;
  signal b1839_flop_next : boolean := false;
  signal b1837_flop_next : boolean := false;
  signal b1835_flop_next : boolean := false;
  signal b1833_flop_next : boolean := false;
  signal b1831_flop_next : boolean := false;
  signal b1829_flop_next : boolean := false;
  signal r1827_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1825_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1823_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1821_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1819_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1817_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1815_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1813_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1811_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1809_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1807_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1805_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1803_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1801_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1799_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1797_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1795_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1792_flop_next : std_logic_vector(0 to 511) := (others => '0');
  signal r1790_flop_next : std_logic_vector(0 to 5) := (others => '0');
  signal r1787_flop_next : std_logic_vector(0 to 5) := (others => '0');
  signal r1783_flop_next : std_logic_vector(0 to 67) := (others => '0');
  signal r1779_flop_next : std_logic_vector(0 to 63) := (others => '0');
  signal r1778_flop_next : std_logic_vector(0 to 64) := (others => '0');
  signal r1776_flop_next : std_logic_vector(0 to 0) := (others => '0');
  signal r1754_flop_next : std_logic_vector(0 to 511) := (others => '0');
  signal b1751_flop_next : boolean := false;
  signal b1749_flop_next : boolean := false;
  signal b1747_flop_next : boolean := false;
  signal b1745_flop_next : boolean := false;
  signal b1743_flop_next : boolean := false;
  signal b1741_flop_next : boolean := false;
  signal b1739_flop_next : boolean := false;
  signal b1737_flop_next : boolean := false;
  signal b1735_flop_next : boolean := false;
  signal b1733_flop_next : boolean := false;
  signal b1731_flop_next : boolean := false;
  signal b1729_flop_next : boolean := false;
  signal b1727_flop_next : boolean := false;
  signal b1725_flop_next : boolean := false;
  signal b1723_flop_next : boolean := false;
  signal b1721_flop_next : boolean := false;
  signal r1719_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1717_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1715_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1713_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1711_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1709_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1707_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1705_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1703_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1701_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1699_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1697_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1695_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1693_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1691_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1689_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal b1686_flop_next : boolean := false;
  signal b1684_flop_next : boolean := false;
  signal r1682_flop_next : std_logic_vector(0 to 511) := (others => '0');
  signal r1680_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1678_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1676_flop_next : std_logic_vector(0 to 511) := (others => '0');
  signal r1670_flop_next : std_logic_vector(0 to 575) := (others => '0');
  signal r1667_flop_next : std_logic_vector(0 to 511) := (others => '0');
  signal r1663_flop_next : std_logic_vector(0 to 255) := (others => '0');
  signal r1659_flop_next : std_logic_vector(0 to 5) := (others => '0');
  signal r1657_flop_next : std_logic_vector(0 to 5) := (others => '0');
  signal b1655_flop_next : boolean := false;
  signal b1653_flop_next : boolean := false;
  signal b1651_flop_next : boolean := false;
  signal r1649_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1647_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal b1645_flop_next : boolean := false;
  signal r1637_flop_next : std_logic_vector(0 to 67) := (others => '0');
  signal r1633_flop_next : std_logic_vector(0 to 63) := (others => '0');
  signal r1632_flop_next : std_logic_vector(0 to 64) := (others => '0');
  signal r1630_flop_next : std_logic_vector(0 to 0) := (others => '0');
  signal r1608_flop_next : std_logic_vector(0 to 511) := (others => '0');
  signal b1605_flop_next : boolean := false;
  signal b1603_flop_next : boolean := false;
  signal b1601_flop_next : boolean := false;
  signal b1599_flop_next : boolean := false;
  signal b1597_flop_next : boolean := false;
  signal b1595_flop_next : boolean := false;
  signal b1593_flop_next : boolean := false;
  signal b1591_flop_next : boolean := false;
  signal b1589_flop_next : boolean := false;
  signal b1587_flop_next : boolean := false;
  signal b1585_flop_next : boolean := false;
  signal b1583_flop_next : boolean := false;
  signal b1581_flop_next : boolean := false;
  signal b1579_flop_next : boolean := false;
  signal b1577_flop_next : boolean := false;
  signal b1575_flop_next : boolean := false;
  signal r1573_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1571_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1569_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1567_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1565_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1563_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1561_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1559_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1557_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1555_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1553_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1551_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1549_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1547_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1545_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1543_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal b1540_flop_next : boolean := false;
  signal b1538_flop_next : boolean := false;
  signal r1536_flop_next : std_logic_vector(0 to 511) := (others => '0');
  signal r1534_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1532_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1530_flop_next : std_logic_vector(0 to 511) := (others => '0');
  signal r1524_flop_next : std_logic_vector(0 to 575) := (others => '0');
  signal r1521_flop_next : std_logic_vector(0 to 511) := (others => '0');
  signal b1519_flop_next : boolean := false;
  signal b1517_flop_next : boolean := false;
  signal b1515_flop_next : boolean := false;
  signal r1513_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1511_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal b1509_flop_next : boolean := false;
  signal r1501_flop_next : std_logic_vector(0 to 67) := (others => '0');
  signal r1497_flop_next : std_logic_vector(0 to 63) := (others => '0');
  signal r1496_flop_next : std_logic_vector(0 to 64) := (others => '0');
  signal r1494_flop_next : std_logic_vector(0 to 0) := (others => '0');
  signal r1472_flop_next : std_logic_vector(0 to 511) := (others => '0');
  signal b1469_flop_next : boolean := false;
  signal b1467_flop_next : boolean := false;
  signal b1465_flop_next : boolean := false;
  signal b1463_flop_next : boolean := false;
  signal b1461_flop_next : boolean := false;
  signal b1459_flop_next : boolean := false;
  signal b1457_flop_next : boolean := false;
  signal b1455_flop_next : boolean := false;
  signal b1453_flop_next : boolean := false;
  signal b1451_flop_next : boolean := false;
  signal b1449_flop_next : boolean := false;
  signal b1447_flop_next : boolean := false;
  signal b1445_flop_next : boolean := false;
  signal b1443_flop_next : boolean := false;
  signal b1441_flop_next : boolean := false;
  signal b1439_flop_next : boolean := false;
  signal r1437_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1435_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1433_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1431_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1429_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1427_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1425_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1423_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1421_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1419_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1417_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1415_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1413_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1411_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1409_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1407_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal b1404_flop_next : boolean := false;
  signal b1402_flop_next : boolean := false;
  signal r1400_flop_next : std_logic_vector(0 to 511) := (others => '0');
  signal r1398_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1396_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1394_flop_next : std_logic_vector(0 to 511) := (others => '0');
  signal r1388_flop_next : std_logic_vector(0 to 575) := (others => '0');
  signal r1385_flop_next : std_logic_vector(0 to 511) := (others => '0');
  signal b1383_flop_next : boolean := false;
  signal b1381_flop_next : boolean := false;
  signal b1379_flop_next : boolean := false;
  signal r1377_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1375_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal b1373_flop_next : boolean := false;
  signal r1365_flop_next : std_logic_vector(0 to 67) := (others => '0');
  signal r1361_flop_next : std_logic_vector(0 to 63) := (others => '0');
  signal r1360_flop_next : std_logic_vector(0 to 64) := (others => '0');
  signal r1358_flop_next : std_logic_vector(0 to 0) := (others => '0');
  signal r1336_flop_next : std_logic_vector(0 to 511) := (others => '0');
  signal b1333_flop_next : boolean := false;
  signal b1331_flop_next : boolean := false;
  signal b1329_flop_next : boolean := false;
  signal b1327_flop_next : boolean := false;
  signal b1325_flop_next : boolean := false;
  signal b1323_flop_next : boolean := false;
  signal b1321_flop_next : boolean := false;
  signal b1319_flop_next : boolean := false;
  signal b1317_flop_next : boolean := false;
  signal b1315_flop_next : boolean := false;
  signal b1313_flop_next : boolean := false;
  signal b1311_flop_next : boolean := false;
  signal b1309_flop_next : boolean := false;
  signal b1307_flop_next : boolean := false;
  signal b1305_flop_next : boolean := false;
  signal b1303_flop_next : boolean := false;
  signal r1301_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1299_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1297_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1295_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1293_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1291_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1289_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1287_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1285_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1283_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1281_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1279_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1277_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1275_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1273_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1271_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal b1268_flop_next : boolean := false;
  signal b1266_flop_next : boolean := false;
  signal r1264_flop_next : std_logic_vector(0 to 511) := (others => '0');
  signal r1262_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1260_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1258_flop_next : std_logic_vector(0 to 511) := (others => '0');
  signal r1252_flop_next : std_logic_vector(0 to 575) := (others => '0');
  signal r1249_flop_next : std_logic_vector(0 to 511) := (others => '0');
  signal b1247_flop_next : boolean := false;
  signal b1245_flop_next : boolean := false;
  signal b1243_flop_next : boolean := false;
  signal r1241_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1239_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal b1237_flop_next : boolean := false;
  signal r1229_flop_next : std_logic_vector(0 to 67) := (others => '0');
  signal r1225_flop_next : std_logic_vector(0 to 63) := (others => '0');
  signal r1224_flop_next : std_logic_vector(0 to 64) := (others => '0');
  signal r1222_flop_next : std_logic_vector(0 to 0) := (others => '0');
  signal r1200_flop_next : std_logic_vector(0 to 511) := (others => '0');
  signal b1197_flop_next : boolean := false;
  signal b1195_flop_next : boolean := false;
  signal b1193_flop_next : boolean := false;
  signal b1191_flop_next : boolean := false;
  signal b1189_flop_next : boolean := false;
  signal b1187_flop_next : boolean := false;
  signal b1185_flop_next : boolean := false;
  signal b1183_flop_next : boolean := false;
  signal b1181_flop_next : boolean := false;
  signal b1179_flop_next : boolean := false;
  signal b1177_flop_next : boolean := false;
  signal b1175_flop_next : boolean := false;
  signal b1173_flop_next : boolean := false;
  signal b1171_flop_next : boolean := false;
  signal b1169_flop_next : boolean := false;
  signal b1167_flop_next : boolean := false;
  signal r1165_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1163_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1161_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1159_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1157_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1155_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1153_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1151_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1149_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1147_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1145_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1143_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1141_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1139_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1137_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1135_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal b1132_flop_next : boolean := false;
  signal b1130_flop_next : boolean := false;
  signal r1128_flop_next : std_logic_vector(0 to 511) := (others => '0');
  signal r1126_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1124_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1122_flop_next : std_logic_vector(0 to 511) := (others => '0');
  signal r1116_flop_next : std_logic_vector(0 to 575) := (others => '0');
  signal r1113_flop_next : std_logic_vector(0 to 511) := (others => '0');
  signal b1111_flop_next : boolean := false;
  signal b1109_flop_next : boolean := false;
  signal b1107_flop_next : boolean := false;
  signal r1105_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1103_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal b1101_flop_next : boolean := false;
  signal r1093_flop_next : std_logic_vector(0 to 67) := (others => '0');
  signal r1089_flop_next : std_logic_vector(0 to 63) := (others => '0');
  signal r1088_flop_next : std_logic_vector(0 to 64) := (others => '0');
  signal r1086_flop_next : std_logic_vector(0 to 0) := (others => '0');
  signal r1064_flop_next : std_logic_vector(0 to 511) := (others => '0');
  signal b1061_flop_next : boolean := false;
  signal b1059_flop_next : boolean := false;
  signal b1057_flop_next : boolean := false;
  signal b1055_flop_next : boolean := false;
  signal b1053_flop_next : boolean := false;
  signal b1051_flop_next : boolean := false;
  signal b1049_flop_next : boolean := false;
  signal b1047_flop_next : boolean := false;
  signal b1045_flop_next : boolean := false;
  signal b1043_flop_next : boolean := false;
  signal b1041_flop_next : boolean := false;
  signal b1039_flop_next : boolean := false;
  signal b1037_flop_next : boolean := false;
  signal b1035_flop_next : boolean := false;
  signal b1033_flop_next : boolean := false;
  signal b1031_flop_next : boolean := false;
  signal r1029_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1027_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1025_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1023_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1021_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1019_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1017_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1015_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1013_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1011_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1009_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1007_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1005_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1003_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1001_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r999_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal b996_flop_next : boolean := false;
  signal b994_flop_next : boolean := false;
  signal r992_flop_next : std_logic_vector(0 to 511) := (others => '0');
  signal r990_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r988_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r986_flop_next : std_logic_vector(0 to 511) := (others => '0');
  signal r980_flop_next : std_logic_vector(0 to 575) := (others => '0');
  signal r977_flop_next : std_logic_vector(0 to 511) := (others => '0');
  signal b975_flop_next : boolean := false;
  signal b973_flop_next : boolean := false;
  signal b971_flop_next : boolean := false;
  signal r969_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r967_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal b965_flop_next : boolean := false;
  signal r957_flop_next : std_logic_vector(0 to 67) := (others => '0');
  signal r953_flop_next : std_logic_vector(0 to 63) := (others => '0');
  signal r952_flop_next : std_logic_vector(0 to 64) := (others => '0');
  signal r950_flop_next : std_logic_vector(0 to 0) := (others => '0');
  signal r928_flop_next : std_logic_vector(0 to 511) := (others => '0');
  signal b925_flop_next : boolean := false;
  signal b923_flop_next : boolean := false;
  signal b921_flop_next : boolean := false;
  signal b919_flop_next : boolean := false;
  signal b917_flop_next : boolean := false;
  signal b915_flop_next : boolean := false;
  signal b913_flop_next : boolean := false;
  signal b911_flop_next : boolean := false;
  signal b909_flop_next : boolean := false;
  signal b907_flop_next : boolean := false;
  signal b905_flop_next : boolean := false;
  signal b903_flop_next : boolean := false;
  signal b901_flop_next : boolean := false;
  signal b899_flop_next : boolean := false;
  signal b897_flop_next : boolean := false;
  signal b895_flop_next : boolean := false;
  signal r893_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r891_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r889_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r887_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r885_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r883_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r881_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r879_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r877_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r875_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r873_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r871_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r869_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r867_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r865_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r863_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal b860_flop_next : boolean := false;
  signal b858_flop_next : boolean := false;
  signal r856_flop_next : std_logic_vector(0 to 511) := (others => '0');
  signal r854_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r852_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r850_flop_next : std_logic_vector(0 to 511) := (others => '0');
  signal r844_flop_next : std_logic_vector(0 to 575) := (others => '0');
  signal r841_flop_next : std_logic_vector(0 to 511) := (others => '0');
  signal b839_flop_next : boolean := false;
  signal b837_flop_next : boolean := false;
  signal b835_flop_next : boolean := false;
  signal r833_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r831_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal b829_flop_next : boolean := false;
  signal r821_flop_next : std_logic_vector(0 to 67) := (others => '0');
  signal r817_flop_next : std_logic_vector(0 to 63) := (others => '0');
  signal r816_flop_next : std_logic_vector(0 to 64) := (others => '0');
  signal r814_flop_next : std_logic_vector(0 to 0) := (others => '0');
  signal r792_flop_next : std_logic_vector(0 to 511) := (others => '0');
  signal b789_flop_next : boolean := false;
  signal b787_flop_next : boolean := false;
  signal b785_flop_next : boolean := false;
  signal b783_flop_next : boolean := false;
  signal b781_flop_next : boolean := false;
  signal b779_flop_next : boolean := false;
  signal b777_flop_next : boolean := false;
  signal b775_flop_next : boolean := false;
  signal b773_flop_next : boolean := false;
  signal b771_flop_next : boolean := false;
  signal b769_flop_next : boolean := false;
  signal b767_flop_next : boolean := false;
  signal b765_flop_next : boolean := false;
  signal b763_flop_next : boolean := false;
  signal b761_flop_next : boolean := false;
  signal b759_flop_next : boolean := false;
  signal r757_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r755_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r753_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r751_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r749_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r747_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r745_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r743_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r741_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r739_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r737_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r735_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r733_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r731_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r729_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r727_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal b724_flop_next : boolean := false;
  signal b722_flop_next : boolean := false;
  signal r720_flop_next : std_logic_vector(0 to 511) := (others => '0');
  signal r718_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r716_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r714_flop_next : std_logic_vector(0 to 511) := (others => '0');
  signal r708_flop_next : std_logic_vector(0 to 575) := (others => '0');
  signal r705_flop_next : std_logic_vector(0 to 511) := (others => '0');
  signal b703_flop_next : boolean := false;
  signal b701_flop_next : boolean := false;
  signal b699_flop_next : boolean := false;
  signal r697_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r695_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal b693_flop_next : boolean := false;
  signal r685_flop_next : std_logic_vector(0 to 67) := (others => '0');
  signal r681_flop_next : std_logic_vector(0 to 63) := (others => '0');
  signal r680_flop_next : std_logic_vector(0 to 64) := (others => '0');
  signal r678_flop_next : std_logic_vector(0 to 0) := (others => '0');
  signal r656_flop_next : std_logic_vector(0 to 511) := (others => '0');
  signal b653_flop_next : boolean := false;
  signal b651_flop_next : boolean := false;
  signal b649_flop_next : boolean := false;
  signal b647_flop_next : boolean := false;
  signal b645_flop_next : boolean := false;
  signal b643_flop_next : boolean := false;
  signal b641_flop_next : boolean := false;
  signal b639_flop_next : boolean := false;
  signal b637_flop_next : boolean := false;
  signal b635_flop_next : boolean := false;
  signal b633_flop_next : boolean := false;
  signal b631_flop_next : boolean := false;
  signal b629_flop_next : boolean := false;
  signal b627_flop_next : boolean := false;
  signal b625_flop_next : boolean := false;
  signal b623_flop_next : boolean := false;
  signal r621_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r619_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r617_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r615_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r613_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r611_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r609_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r607_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r605_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r603_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r601_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r599_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r597_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r595_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r593_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r591_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal b588_flop_next : boolean := false;
  signal b586_flop_next : boolean := false;
  signal r584_flop_next : std_logic_vector(0 to 511) := (others => '0');
  signal r582_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r580_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r578_flop_next : std_logic_vector(0 to 511) := (others => '0');
  signal r572_flop_next : std_logic_vector(0 to 575) := (others => '0');
  signal r569_flop_next : std_logic_vector(0 to 511) := (others => '0');
  signal r566_flop_next : std_logic_vector(0 to 255) := (others => '0');
  signal b26_flop_next : boolean := false;
  signal b24_flop_next : boolean := false;
  signal b22_flop_next : boolean := false;
  signal r20_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r18_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal b16_flop_next : boolean := false;
  signal r12_flop_next : std_logic_vector(0 to 67) := (others => '0');
  signal r10_flop_next : std_logic_vector(0 to 67) := (others => '0');
  signal r6_flop_next : std_logic_vector(0 to 63) := (others => '0');
  signal r5_flop_next : std_logic_vector(0 to 64) := (others => '0');
  signal r3_flop_next : std_logic_vector(0 to 0) := (others => '0');
  signal statevar0_flop_next : std_logic_vector(0 to 255) := (others => '0');
  signal statevar1_flop_next : std_logic_vector(0 to 511) := (others => '0');
  signal statevar2_flop_next : std_logic_vector(0 to 255) := (others => '0');
  signal statevar3_flop_next : std_logic_vector(0 to 5) := (others => '0');
begin
  -- Logic loop process.
  process (control_flop,input_flop,goto_L7851_flop,goto_L7844_flop,goto_L7806_flop,goto_L7767_flop,goto_L7728_flop,goto_L7570_flop,goto_L7690_flop,goto_L7575_flop,goto_L1784_flop,goto_L1785_flop,goto_L1638_flop,goto_L1502_flop,goto_L1366_flop,goto_L1230_flop,goto_L1094_flop,goto_L958_flop,goto_L822_flop,goto_L686_flop,goto_L11_flop,goto_L13_flop,goto_L690_flop,goto_L826_flop,goto_L962_flop,goto_L1098_flop,goto_L1234_flop,goto_L1370_flop,goto_L1506_flop,goto_L1642_flop,goto_L7693_flop,goto_L7732_flop,goto_L7771_flop,goto_L7810_flop,goto_L7777_flop,goto_L7738_flop,goto_L7699_flop,goto_L1658_flop,goto_L1522_flop,goto_L1386_flop,goto_L1250_flop,goto_L1114_flop,goto_L978_flop,goto_L842_flop,goto_L706_flop,goto_L567_flop,goto_L0_flop,goto_L7852_flop,r7843_flop,r7840_flop,r7817_flop,r7814_flop,r7805_flop,r7802_flop,r7779_flop,r7776_flop,b7774_flop,r7766_flop,r7763_flop,r7740_flop,r7737_flop,b7735_flop,r7727_flop,r7724_flop,r7701_flop,r7698_flop,b7696_flop,r7679_flop,r7675_flop,r7671_flop,r7667_flop,r7663_flop,r7659_flop,r7655_flop,r7651_flop,r7647_flop,b7644_flop,b7642_flop,b7640_flop,b7638_flop,b7636_flop,b7634_flop,b7632_flop,b7630_flop,r7628_flop,r7626_flop,r7624_flop,r7622_flop,r7620_flop,r7618_flop,r7616_flop,r7614_flop,r7610_flop,b7608_flop,b7606_flop,b7604_flop,b7602_flop,b7600_flop,b7598_flop,b7596_flop,b7594_flop,r7592_flop,r7590_flop,r7588_flop,r7586_flop,r7584_flop,r7582_flop,r7580_flop,r7578_flop,r7574_flop,b7572_flop,r7569_flop,r7565_flop,r7564_flop,r7562_flop,r7558_flop,r7300_flop,r7296_flop,r7292_flop,r2874_flop,r2376_flop,r2375_flop,r2374_flop,r2371_flop,r2365_flop,r1862_flop,b1859_flop,b1857_flop,b1855_flop,b1853_flop,b1851_flop,b1849_flop,b1847_flop,b1845_flop,b1843_flop,b1841_flop,b1839_flop,b1837_flop,b1835_flop,b1833_flop,b1831_flop,b1829_flop,r1827_flop,r1825_flop,r1823_flop,r1821_flop,r1819_flop,r1817_flop,r1815_flop,r1813_flop,r1811_flop,r1809_flop,r1807_flop,r1805_flop,r1803_flop,r1801_flop,r1799_flop,r1797_flop,r1795_flop,r1792_flop,r1790_flop,r1787_flop,r1783_flop,r1779_flop,r1778_flop,r1776_flop,r1754_flop,b1751_flop,b1749_flop,b1747_flop,b1745_flop,b1743_flop,b1741_flop,b1739_flop,b1737_flop,b1735_flop,b1733_flop,b1731_flop,b1729_flop,b1727_flop,b1725_flop,b1723_flop,b1721_flop,r1719_flop,r1717_flop,r1715_flop,r1713_flop,r1711_flop,r1709_flop,r1707_flop,r1705_flop,r1703_flop,r1701_flop,r1699_flop,r1697_flop,r1695_flop,r1693_flop,r1691_flop,r1689_flop,b1686_flop,b1684_flop,r1682_flop,r1680_flop,r1678_flop,r1676_flop,r1670_flop,r1667_flop,r1663_flop,r1659_flop,r1657_flop,b1655_flop,b1653_flop,b1651_flop,r1649_flop,r1647_flop,b1645_flop,r1637_flop,r1633_flop,r1632_flop,r1630_flop,r1608_flop,b1605_flop,b1603_flop,b1601_flop,b1599_flop,b1597_flop,b1595_flop,b1593_flop,b1591_flop,b1589_flop,b1587_flop,b1585_flop,b1583_flop,b1581_flop,b1579_flop,b1577_flop,b1575_flop,r1573_flop,r1571_flop,r1569_flop,r1567_flop,r1565_flop,r1563_flop,r1561_flop,r1559_flop,r1557_flop,r1555_flop,r1553_flop,r1551_flop,r1549_flop,r1547_flop,r1545_flop,r1543_flop,b1540_flop,b1538_flop,r1536_flop,r1534_flop,r1532_flop,r1530_flop,r1524_flop,r1521_flop,b1519_flop,b1517_flop,b1515_flop,r1513_flop,r1511_flop,b1509_flop,r1501_flop,r1497_flop,r1496_flop,r1494_flop,r1472_flop,b1469_flop,b1467_flop,b1465_flop,b1463_flop,b1461_flop,b1459_flop,b1457_flop,b1455_flop,b1453_flop,b1451_flop,b1449_flop,b1447_flop,b1445_flop,b1443_flop,b1441_flop,b1439_flop,r1437_flop,r1435_flop,r1433_flop,r1431_flop,r1429_flop,r1427_flop,r1425_flop,r1423_flop,r1421_flop,r1419_flop,r1417_flop,r1415_flop,r1413_flop,r1411_flop,r1409_flop,r1407_flop,b1404_flop,b1402_flop,r1400_flop,r1398_flop,r1396_flop,r1394_flop,r1388_flop,r1385_flop,b1383_flop,b1381_flop,b1379_flop,r1377_flop,r1375_flop,b1373_flop,r1365_flop,r1361_flop,r1360_flop,r1358_flop,r1336_flop,b1333_flop,b1331_flop,b1329_flop,b1327_flop,b1325_flop,b1323_flop,b1321_flop,b1319_flop,b1317_flop,b1315_flop,b1313_flop,b1311_flop,b1309_flop,b1307_flop,b1305_flop,b1303_flop,r1301_flop,r1299_flop,r1297_flop,r1295_flop,r1293_flop,r1291_flop,r1289_flop,r1287_flop,r1285_flop,r1283_flop,r1281_flop,r1279_flop,r1277_flop,r1275_flop,r1273_flop,r1271_flop,b1268_flop,b1266_flop,r1264_flop,r1262_flop,r1260_flop,r1258_flop,r1252_flop,r1249_flop,b1247_flop,b1245_flop,b1243_flop,r1241_flop,r1239_flop,b1237_flop,r1229_flop,r1225_flop,r1224_flop,r1222_flop,r1200_flop,b1197_flop,b1195_flop,b1193_flop,b1191_flop,b1189_flop,b1187_flop,b1185_flop,b1183_flop,b1181_flop,b1179_flop,b1177_flop,b1175_flop,b1173_flop,b1171_flop,b1169_flop,b1167_flop,r1165_flop,r1163_flop,r1161_flop,r1159_flop,r1157_flop,r1155_flop,r1153_flop,r1151_flop,r1149_flop,r1147_flop,r1145_flop,r1143_flop,r1141_flop,r1139_flop,r1137_flop,r1135_flop,b1132_flop,b1130_flop,r1128_flop,r1126_flop,r1124_flop,r1122_flop,r1116_flop,r1113_flop,b1111_flop,b1109_flop,b1107_flop,r1105_flop,r1103_flop,b1101_flop,r1093_flop,r1089_flop,r1088_flop,r1086_flop,r1064_flop,b1061_flop,b1059_flop,b1057_flop,b1055_flop,b1053_flop,b1051_flop,b1049_flop,b1047_flop,b1045_flop,b1043_flop,b1041_flop,b1039_flop,b1037_flop,b1035_flop,b1033_flop,b1031_flop,r1029_flop,r1027_flop,r1025_flop,r1023_flop,r1021_flop,r1019_flop,r1017_flop,r1015_flop,r1013_flop,r1011_flop,r1009_flop,r1007_flop,r1005_flop,r1003_flop,r1001_flop,r999_flop,b996_flop,b994_flop,r992_flop,r990_flop,r988_flop,r986_flop,r980_flop,r977_flop,b975_flop,b973_flop,b971_flop,r969_flop,r967_flop,b965_flop,r957_flop,r953_flop,r952_flop,r950_flop,r928_flop,b925_flop,b923_flop,b921_flop,b919_flop,b917_flop,b915_flop,b913_flop,b911_flop,b909_flop,b907_flop,b905_flop,b903_flop,b901_flop,b899_flop,b897_flop,b895_flop,r893_flop,r891_flop,r889_flop,r887_flop,r885_flop,r883_flop,r881_flop,r879_flop,r877_flop,r875_flop,r873_flop,r871_flop,r869_flop,r867_flop,r865_flop,r863_flop,b860_flop,b858_flop,r856_flop,r854_flop,r852_flop,r850_flop,r844_flop,r841_flop,b839_flop,b837_flop,b835_flop,r833_flop,r831_flop,b829_flop,r821_flop,r817_flop,r816_flop,r814_flop,r792_flop,b789_flop,b787_flop,b785_flop,b783_flop,b781_flop,b779_flop,b777_flop,b775_flop,b773_flop,b771_flop,b769_flop,b767_flop,b765_flop,b763_flop,b761_flop,b759_flop,r757_flop,r755_flop,r753_flop,r751_flop,r749_flop,r747_flop,r745_flop,r743_flop,r741_flop,r739_flop,r737_flop,r735_flop,r733_flop,r731_flop,r729_flop,r727_flop,b724_flop,b722_flop,r720_flop,r718_flop,r716_flop,r714_flop,r708_flop,r705_flop,b703_flop,b701_flop,b699_flop,r697_flop,r695_flop,b693_flop,r685_flop,r681_flop,r680_flop,r678_flop,r656_flop,b653_flop,b651_flop,b649_flop,b647_flop,b645_flop,b643_flop,b641_flop,b639_flop,b637_flop,b635_flop,b633_flop,b631_flop,b629_flop,b627_flop,b625_flop,b623_flop,r621_flop,r619_flop,r617_flop,r615_flop,r613_flop,r611_flop,r609_flop,r607_flop,r605_flop,r603_flop,r601_flop,r599_flop,r597_flop,r595_flop,r593_flop,r591_flop,b588_flop,b586_flop,r584_flop,r582_flop,r580_flop,r578_flop,r572_flop,r569_flop,r566_flop,b26_flop,b24_flop,b22_flop,r20_flop,r18_flop,b16_flop,r12_flop,r10_flop,r6_flop,r5_flop,r3_flop,statevar0_flop,statevar1_flop,statevar2_flop,statevar3_flop)
    variable control : control_state;
    variable input_tmp : std_logic_vector(0 to 67);
    variable goto_L7851 : boolean := false;
    variable goto_L7844 : boolean := false;
    variable goto_L7806 : boolean := false;
    variable goto_L7767 : boolean := false;
    variable goto_L7728 : boolean := false;
    variable goto_L7570 : boolean := false;
    variable goto_L7690 : boolean := false;
    variable goto_L7575 : boolean := false;
    variable goto_L1784 : boolean := false;
    variable goto_L1785 : boolean := false;
    variable goto_L1638 : boolean := false;
    variable goto_L1502 : boolean := false;
    variable goto_L1366 : boolean := false;
    variable goto_L1230 : boolean := false;
    variable goto_L1094 : boolean := false;
    variable goto_L958 : boolean := false;
    variable goto_L822 : boolean := false;
    variable goto_L686 : boolean := false;
    variable goto_L11 : boolean := false;
    variable goto_L13 : boolean := false;
    variable goto_L690 : boolean := false;
    variable goto_L826 : boolean := false;
    variable goto_L962 : boolean := false;
    variable goto_L1098 : boolean := false;
    variable goto_L1234 : boolean := false;
    variable goto_L1370 : boolean := false;
    variable goto_L1506 : boolean := false;
    variable goto_L1642 : boolean := false;
    variable goto_L7693 : boolean := false;
    variable goto_L7732 : boolean := false;
    variable goto_L7771 : boolean := false;
    variable goto_L7810 : boolean := false;
    variable goto_L7777 : boolean := false;
    variable goto_L7738 : boolean := false;
    variable goto_L7699 : boolean := false;
    variable goto_L1658 : boolean := false;
    variable goto_L1522 : boolean := false;
    variable goto_L1386 : boolean := false;
    variable goto_L1250 : boolean := false;
    variable goto_L1114 : boolean := false;
    variable goto_L978 : boolean := false;
    variable goto_L842 : boolean := false;
    variable goto_L706 : boolean := false;
    variable goto_L567 : boolean := false;
    variable goto_L0 : boolean := false;
    variable goto_L7852 : boolean := false;
    variable r7843 : std_logic_vector(0 to 67) := (others => '0');
    variable r7840 : std_logic_vector(0 to 64) := (others => '0');
    variable r7817 : std_logic_vector(0 to 255) := (others => '0');
    variable r7814 : std_logic_vector(0 to 255) := (others => '0');
    variable r7805 : std_logic_vector(0 to 67) := (others => '0');
    variable r7802 : std_logic_vector(0 to 64) := (others => '0');
    variable r7779 : std_logic_vector(0 to 255) := (others => '0');
    variable r7776 : std_logic_vector(0 to 255) := (others => '0');
    variable b7774 : boolean := false;
    variable r7766 : std_logic_vector(0 to 67) := (others => '0');
    variable r7763 : std_logic_vector(0 to 64) := (others => '0');
    variable r7740 : std_logic_vector(0 to 255) := (others => '0');
    variable r7737 : std_logic_vector(0 to 255) := (others => '0');
    variable b7735 : boolean := false;
    variable r7727 : std_logic_vector(0 to 67) := (others => '0');
    variable r7724 : std_logic_vector(0 to 64) := (others => '0');
    variable r7701 : std_logic_vector(0 to 255) := (others => '0');
    variable r7698 : std_logic_vector(0 to 255) := (others => '0');
    variable b7696 : boolean := false;
    variable r7679 : std_logic_vector(0 to 31) := (others => '0');
    variable r7675 : std_logic_vector(0 to 31) := (others => '0');
    variable r7671 : std_logic_vector(0 to 31) := (others => '0');
    variable r7667 : std_logic_vector(0 to 31) := (others => '0');
    variable r7663 : std_logic_vector(0 to 31) := (others => '0');
    variable r7659 : std_logic_vector(0 to 31) := (others => '0');
    variable r7655 : std_logic_vector(0 to 31) := (others => '0');
    variable r7651 : std_logic_vector(0 to 31) := (others => '0');
    variable r7647 : std_logic_vector(0 to 255) := (others => '0');
    variable b7644 : boolean := false;
    variable b7642 : boolean := false;
    variable b7640 : boolean := false;
    variable b7638 : boolean := false;
    variable b7636 : boolean := false;
    variable b7634 : boolean := false;
    variable b7632 : boolean := false;
    variable b7630 : boolean := false;
    variable r7628 : std_logic_vector(0 to 31) := (others => '0');
    variable r7626 : std_logic_vector(0 to 31) := (others => '0');
    variable r7624 : std_logic_vector(0 to 31) := (others => '0');
    variable r7622 : std_logic_vector(0 to 31) := (others => '0');
    variable r7620 : std_logic_vector(0 to 31) := (others => '0');
    variable r7618 : std_logic_vector(0 to 31) := (others => '0');
    variable r7616 : std_logic_vector(0 to 31) := (others => '0');
    variable r7614 : std_logic_vector(0 to 31) := (others => '0');
    variable r7610 : std_logic_vector(0 to 255) := (others => '0');
    variable b7608 : boolean := false;
    variable b7606 : boolean := false;
    variable b7604 : boolean := false;
    variable b7602 : boolean := false;
    variable b7600 : boolean := false;
    variable b7598 : boolean := false;
    variable b7596 : boolean := false;
    variable b7594 : boolean := false;
    variable r7592 : std_logic_vector(0 to 31) := (others => '0');
    variable r7590 : std_logic_vector(0 to 31) := (others => '0');
    variable r7588 : std_logic_vector(0 to 31) := (others => '0');
    variable r7586 : std_logic_vector(0 to 31) := (others => '0');
    variable r7584 : std_logic_vector(0 to 31) := (others => '0');
    variable r7582 : std_logic_vector(0 to 31) := (others => '0');
    variable r7580 : std_logic_vector(0 to 31) := (others => '0');
    variable r7578 : std_logic_vector(0 to 31) := (others => '0');
    variable r7574 : std_logic_vector(0 to 255) := (others => '0');
    variable b7572 : boolean := false;
    variable r7569 : std_logic_vector(0 to 67) := (others => '0');
    variable r7565 : std_logic_vector(0 to 63) := (others => '0');
    variable r7564 : std_logic_vector(0 to 64) := (others => '0');
    variable r7562 : std_logic_vector(0 to 0) := (others => '0');
    variable r7558 : std_logic_vector(0 to 5) := (others => '0');
    variable r7300 : std_logic_vector(0 to 5) := (others => '0');
    variable r7296 : std_logic_vector(0 to 255) := (others => '0');
    variable r7292 : std_logic_vector(0 to 31) := (others => '0');
    variable r2874 : std_logic_vector(0 to 5) := (others => '0');
    variable r2376 : std_logic_vector(0 to 255) := (others => '0');
    variable r2375 : std_logic_vector(0 to 31) := (others => '0');
    variable r2374 : std_logic_vector(0 to 31) := (others => '0');
    variable r2371 : std_logic_vector(0 to 255) := (others => '0');
    variable r2365 : std_logic_vector(0 to 511) := (others => '0');
    variable r1862 : std_logic_vector(0 to 511) := (others => '0');
    variable b1859 : boolean := false;
    variable b1857 : boolean := false;
    variable b1855 : boolean := false;
    variable b1853 : boolean := false;
    variable b1851 : boolean := false;
    variable b1849 : boolean := false;
    variable b1847 : boolean := false;
    variable b1845 : boolean := false;
    variable b1843 : boolean := false;
    variable b1841 : boolean := false;
    variable b1839 : boolean := false;
    variable b1837 : boolean := false;
    variable b1835 : boolean := false;
    variable b1833 : boolean := false;
    variable b1831 : boolean := false;
    variable b1829 : boolean := false;
    variable r1827 : std_logic_vector(0 to 31) := (others => '0');
    variable r1825 : std_logic_vector(0 to 31) := (others => '0');
    variable r1823 : std_logic_vector(0 to 31) := (others => '0');
    variable r1821 : std_logic_vector(0 to 31) := (others => '0');
    variable r1819 : std_logic_vector(0 to 31) := (others => '0');
    variable r1817 : std_logic_vector(0 to 31) := (others => '0');
    variable r1815 : std_logic_vector(0 to 31) := (others => '0');
    variable r1813 : std_logic_vector(0 to 31) := (others => '0');
    variable r1811 : std_logic_vector(0 to 31) := (others => '0');
    variable r1809 : std_logic_vector(0 to 31) := (others => '0');
    variable r1807 : std_logic_vector(0 to 31) := (others => '0');
    variable r1805 : std_logic_vector(0 to 31) := (others => '0');
    variable r1803 : std_logic_vector(0 to 31) := (others => '0');
    variable r1801 : std_logic_vector(0 to 31) := (others => '0');
    variable r1799 : std_logic_vector(0 to 31) := (others => '0');
    variable r1797 : std_logic_vector(0 to 31) := (others => '0');
    variable r1795 : std_logic_vector(0 to 31) := (others => '0');
    variable r1792 : std_logic_vector(0 to 511) := (others => '0');
    variable r1790 : std_logic_vector(0 to 5) := (others => '0');
    variable r1787 : std_logic_vector(0 to 5) := (others => '0');
    variable r1783 : std_logic_vector(0 to 67) := (others => '0');
    variable r1779 : std_logic_vector(0 to 63) := (others => '0');
    variable r1778 : std_logic_vector(0 to 64) := (others => '0');
    variable r1776 : std_logic_vector(0 to 0) := (others => '0');
    variable r1754 : std_logic_vector(0 to 511) := (others => '0');
    variable b1751 : boolean := false;
    variable b1749 : boolean := false;
    variable b1747 : boolean := false;
    variable b1745 : boolean := false;
    variable b1743 : boolean := false;
    variable b1741 : boolean := false;
    variable b1739 : boolean := false;
    variable b1737 : boolean := false;
    variable b1735 : boolean := false;
    variable b1733 : boolean := false;
    variable b1731 : boolean := false;
    variable b1729 : boolean := false;
    variable b1727 : boolean := false;
    variable b1725 : boolean := false;
    variable b1723 : boolean := false;
    variable b1721 : boolean := false;
    variable r1719 : std_logic_vector(0 to 31) := (others => '0');
    variable r1717 : std_logic_vector(0 to 31) := (others => '0');
    variable r1715 : std_logic_vector(0 to 31) := (others => '0');
    variable r1713 : std_logic_vector(0 to 31) := (others => '0');
    variable r1711 : std_logic_vector(0 to 31) := (others => '0');
    variable r1709 : std_logic_vector(0 to 31) := (others => '0');
    variable r1707 : std_logic_vector(0 to 31) := (others => '0');
    variable r1705 : std_logic_vector(0 to 31) := (others => '0');
    variable r1703 : std_logic_vector(0 to 31) := (others => '0');
    variable r1701 : std_logic_vector(0 to 31) := (others => '0');
    variable r1699 : std_logic_vector(0 to 31) := (others => '0');
    variable r1697 : std_logic_vector(0 to 31) := (others => '0');
    variable r1695 : std_logic_vector(0 to 31) := (others => '0');
    variable r1693 : std_logic_vector(0 to 31) := (others => '0');
    variable r1691 : std_logic_vector(0 to 31) := (others => '0');
    variable r1689 : std_logic_vector(0 to 31) := (others => '0');
    variable b1686 : boolean := false;
    variable b1684 : boolean := false;
    variable r1682 : std_logic_vector(0 to 511) := (others => '0');
    variable r1680 : std_logic_vector(0 to 31) := (others => '0');
    variable r1678 : std_logic_vector(0 to 31) := (others => '0');
    variable r1676 : std_logic_vector(0 to 511) := (others => '0');
    variable r1670 : std_logic_vector(0 to 575) := (others => '0');
    variable r1667 : std_logic_vector(0 to 511) := (others => '0');
    variable r1663 : std_logic_vector(0 to 255) := (others => '0');
    variable r1659 : std_logic_vector(0 to 5) := (others => '0');
    variable r1657 : std_logic_vector(0 to 5) := (others => '0');
    variable b1655 : boolean := false;
    variable b1653 : boolean := false;
    variable b1651 : boolean := false;
    variable r1649 : std_logic_vector(0 to 31) := (others => '0');
    variable r1647 : std_logic_vector(0 to 31) := (others => '0');
    variable b1645 : boolean := false;
    variable r1637 : std_logic_vector(0 to 67) := (others => '0');
    variable r1633 : std_logic_vector(0 to 63) := (others => '0');
    variable r1632 : std_logic_vector(0 to 64) := (others => '0');
    variable r1630 : std_logic_vector(0 to 0) := (others => '0');
    variable r1608 : std_logic_vector(0 to 511) := (others => '0');
    variable b1605 : boolean := false;
    variable b1603 : boolean := false;
    variable b1601 : boolean := false;
    variable b1599 : boolean := false;
    variable b1597 : boolean := false;
    variable b1595 : boolean := false;
    variable b1593 : boolean := false;
    variable b1591 : boolean := false;
    variable b1589 : boolean := false;
    variable b1587 : boolean := false;
    variable b1585 : boolean := false;
    variable b1583 : boolean := false;
    variable b1581 : boolean := false;
    variable b1579 : boolean := false;
    variable b1577 : boolean := false;
    variable b1575 : boolean := false;
    variable r1573 : std_logic_vector(0 to 31) := (others => '0');
    variable r1571 : std_logic_vector(0 to 31) := (others => '0');
    variable r1569 : std_logic_vector(0 to 31) := (others => '0');
    variable r1567 : std_logic_vector(0 to 31) := (others => '0');
    variable r1565 : std_logic_vector(0 to 31) := (others => '0');
    variable r1563 : std_logic_vector(0 to 31) := (others => '0');
    variable r1561 : std_logic_vector(0 to 31) := (others => '0');
    variable r1559 : std_logic_vector(0 to 31) := (others => '0');
    variable r1557 : std_logic_vector(0 to 31) := (others => '0');
    variable r1555 : std_logic_vector(0 to 31) := (others => '0');
    variable r1553 : std_logic_vector(0 to 31) := (others => '0');
    variable r1551 : std_logic_vector(0 to 31) := (others => '0');
    variable r1549 : std_logic_vector(0 to 31) := (others => '0');
    variable r1547 : std_logic_vector(0 to 31) := (others => '0');
    variable r1545 : std_logic_vector(0 to 31) := (others => '0');
    variable r1543 : std_logic_vector(0 to 31) := (others => '0');
    variable b1540 : boolean := false;
    variable b1538 : boolean := false;
    variable r1536 : std_logic_vector(0 to 511) := (others => '0');
    variable r1534 : std_logic_vector(0 to 31) := (others => '0');
    variable r1532 : std_logic_vector(0 to 31) := (others => '0');
    variable r1530 : std_logic_vector(0 to 511) := (others => '0');
    variable r1524 : std_logic_vector(0 to 575) := (others => '0');
    variable r1521 : std_logic_vector(0 to 511) := (others => '0');
    variable b1519 : boolean := false;
    variable b1517 : boolean := false;
    variable b1515 : boolean := false;
    variable r1513 : std_logic_vector(0 to 31) := (others => '0');
    variable r1511 : std_logic_vector(0 to 31) := (others => '0');
    variable b1509 : boolean := false;
    variable r1501 : std_logic_vector(0 to 67) := (others => '0');
    variable r1497 : std_logic_vector(0 to 63) := (others => '0');
    variable r1496 : std_logic_vector(0 to 64) := (others => '0');
    variable r1494 : std_logic_vector(0 to 0) := (others => '0');
    variable r1472 : std_logic_vector(0 to 511) := (others => '0');
    variable b1469 : boolean := false;
    variable b1467 : boolean := false;
    variable b1465 : boolean := false;
    variable b1463 : boolean := false;
    variable b1461 : boolean := false;
    variable b1459 : boolean := false;
    variable b1457 : boolean := false;
    variable b1455 : boolean := false;
    variable b1453 : boolean := false;
    variable b1451 : boolean := false;
    variable b1449 : boolean := false;
    variable b1447 : boolean := false;
    variable b1445 : boolean := false;
    variable b1443 : boolean := false;
    variable b1441 : boolean := false;
    variable b1439 : boolean := false;
    variable r1437 : std_logic_vector(0 to 31) := (others => '0');
    variable r1435 : std_logic_vector(0 to 31) := (others => '0');
    variable r1433 : std_logic_vector(0 to 31) := (others => '0');
    variable r1431 : std_logic_vector(0 to 31) := (others => '0');
    variable r1429 : std_logic_vector(0 to 31) := (others => '0');
    variable r1427 : std_logic_vector(0 to 31) := (others => '0');
    variable r1425 : std_logic_vector(0 to 31) := (others => '0');
    variable r1423 : std_logic_vector(0 to 31) := (others => '0');
    variable r1421 : std_logic_vector(0 to 31) := (others => '0');
    variable r1419 : std_logic_vector(0 to 31) := (others => '0');
    variable r1417 : std_logic_vector(0 to 31) := (others => '0');
    variable r1415 : std_logic_vector(0 to 31) := (others => '0');
    variable r1413 : std_logic_vector(0 to 31) := (others => '0');
    variable r1411 : std_logic_vector(0 to 31) := (others => '0');
    variable r1409 : std_logic_vector(0 to 31) := (others => '0');
    variable r1407 : std_logic_vector(0 to 31) := (others => '0');
    variable b1404 : boolean := false;
    variable b1402 : boolean := false;
    variable r1400 : std_logic_vector(0 to 511) := (others => '0');
    variable r1398 : std_logic_vector(0 to 31) := (others => '0');
    variable r1396 : std_logic_vector(0 to 31) := (others => '0');
    variable r1394 : std_logic_vector(0 to 511) := (others => '0');
    variable r1388 : std_logic_vector(0 to 575) := (others => '0');
    variable r1385 : std_logic_vector(0 to 511) := (others => '0');
    variable b1383 : boolean := false;
    variable b1381 : boolean := false;
    variable b1379 : boolean := false;
    variable r1377 : std_logic_vector(0 to 31) := (others => '0');
    variable r1375 : std_logic_vector(0 to 31) := (others => '0');
    variable b1373 : boolean := false;
    variable r1365 : std_logic_vector(0 to 67) := (others => '0');
    variable r1361 : std_logic_vector(0 to 63) := (others => '0');
    variable r1360 : std_logic_vector(0 to 64) := (others => '0');
    variable r1358 : std_logic_vector(0 to 0) := (others => '0');
    variable r1336 : std_logic_vector(0 to 511) := (others => '0');
    variable b1333 : boolean := false;
    variable b1331 : boolean := false;
    variable b1329 : boolean := false;
    variable b1327 : boolean := false;
    variable b1325 : boolean := false;
    variable b1323 : boolean := false;
    variable b1321 : boolean := false;
    variable b1319 : boolean := false;
    variable b1317 : boolean := false;
    variable b1315 : boolean := false;
    variable b1313 : boolean := false;
    variable b1311 : boolean := false;
    variable b1309 : boolean := false;
    variable b1307 : boolean := false;
    variable b1305 : boolean := false;
    variable b1303 : boolean := false;
    variable r1301 : std_logic_vector(0 to 31) := (others => '0');
    variable r1299 : std_logic_vector(0 to 31) := (others => '0');
    variable r1297 : std_logic_vector(0 to 31) := (others => '0');
    variable r1295 : std_logic_vector(0 to 31) := (others => '0');
    variable r1293 : std_logic_vector(0 to 31) := (others => '0');
    variable r1291 : std_logic_vector(0 to 31) := (others => '0');
    variable r1289 : std_logic_vector(0 to 31) := (others => '0');
    variable r1287 : std_logic_vector(0 to 31) := (others => '0');
    variable r1285 : std_logic_vector(0 to 31) := (others => '0');
    variable r1283 : std_logic_vector(0 to 31) := (others => '0');
    variable r1281 : std_logic_vector(0 to 31) := (others => '0');
    variable r1279 : std_logic_vector(0 to 31) := (others => '0');
    variable r1277 : std_logic_vector(0 to 31) := (others => '0');
    variable r1275 : std_logic_vector(0 to 31) := (others => '0');
    variable r1273 : std_logic_vector(0 to 31) := (others => '0');
    variable r1271 : std_logic_vector(0 to 31) := (others => '0');
    variable b1268 : boolean := false;
    variable b1266 : boolean := false;
    variable r1264 : std_logic_vector(0 to 511) := (others => '0');
    variable r1262 : std_logic_vector(0 to 31) := (others => '0');
    variable r1260 : std_logic_vector(0 to 31) := (others => '0');
    variable r1258 : std_logic_vector(0 to 511) := (others => '0');
    variable r1252 : std_logic_vector(0 to 575) := (others => '0');
    variable r1249 : std_logic_vector(0 to 511) := (others => '0');
    variable b1247 : boolean := false;
    variable b1245 : boolean := false;
    variable b1243 : boolean := false;
    variable r1241 : std_logic_vector(0 to 31) := (others => '0');
    variable r1239 : std_logic_vector(0 to 31) := (others => '0');
    variable b1237 : boolean := false;
    variable r1229 : std_logic_vector(0 to 67) := (others => '0');
    variable r1225 : std_logic_vector(0 to 63) := (others => '0');
    variable r1224 : std_logic_vector(0 to 64) := (others => '0');
    variable r1222 : std_logic_vector(0 to 0) := (others => '0');
    variable r1200 : std_logic_vector(0 to 511) := (others => '0');
    variable b1197 : boolean := false;
    variable b1195 : boolean := false;
    variable b1193 : boolean := false;
    variable b1191 : boolean := false;
    variable b1189 : boolean := false;
    variable b1187 : boolean := false;
    variable b1185 : boolean := false;
    variable b1183 : boolean := false;
    variable b1181 : boolean := false;
    variable b1179 : boolean := false;
    variable b1177 : boolean := false;
    variable b1175 : boolean := false;
    variable b1173 : boolean := false;
    variable b1171 : boolean := false;
    variable b1169 : boolean := false;
    variable b1167 : boolean := false;
    variable r1165 : std_logic_vector(0 to 31) := (others => '0');
    variable r1163 : std_logic_vector(0 to 31) := (others => '0');
    variable r1161 : std_logic_vector(0 to 31) := (others => '0');
    variable r1159 : std_logic_vector(0 to 31) := (others => '0');
    variable r1157 : std_logic_vector(0 to 31) := (others => '0');
    variable r1155 : std_logic_vector(0 to 31) := (others => '0');
    variable r1153 : std_logic_vector(0 to 31) := (others => '0');
    variable r1151 : std_logic_vector(0 to 31) := (others => '0');
    variable r1149 : std_logic_vector(0 to 31) := (others => '0');
    variable r1147 : std_logic_vector(0 to 31) := (others => '0');
    variable r1145 : std_logic_vector(0 to 31) := (others => '0');
    variable r1143 : std_logic_vector(0 to 31) := (others => '0');
    variable r1141 : std_logic_vector(0 to 31) := (others => '0');
    variable r1139 : std_logic_vector(0 to 31) := (others => '0');
    variable r1137 : std_logic_vector(0 to 31) := (others => '0');
    variable r1135 : std_logic_vector(0 to 31) := (others => '0');
    variable b1132 : boolean := false;
    variable b1130 : boolean := false;
    variable r1128 : std_logic_vector(0 to 511) := (others => '0');
    variable r1126 : std_logic_vector(0 to 31) := (others => '0');
    variable r1124 : std_logic_vector(0 to 31) := (others => '0');
    variable r1122 : std_logic_vector(0 to 511) := (others => '0');
    variable r1116 : std_logic_vector(0 to 575) := (others => '0');
    variable r1113 : std_logic_vector(0 to 511) := (others => '0');
    variable b1111 : boolean := false;
    variable b1109 : boolean := false;
    variable b1107 : boolean := false;
    variable r1105 : std_logic_vector(0 to 31) := (others => '0');
    variable r1103 : std_logic_vector(0 to 31) := (others => '0');
    variable b1101 : boolean := false;
    variable r1093 : std_logic_vector(0 to 67) := (others => '0');
    variable r1089 : std_logic_vector(0 to 63) := (others => '0');
    variable r1088 : std_logic_vector(0 to 64) := (others => '0');
    variable r1086 : std_logic_vector(0 to 0) := (others => '0');
    variable r1064 : std_logic_vector(0 to 511) := (others => '0');
    variable b1061 : boolean := false;
    variable b1059 : boolean := false;
    variable b1057 : boolean := false;
    variable b1055 : boolean := false;
    variable b1053 : boolean := false;
    variable b1051 : boolean := false;
    variable b1049 : boolean := false;
    variable b1047 : boolean := false;
    variable b1045 : boolean := false;
    variable b1043 : boolean := false;
    variable b1041 : boolean := false;
    variable b1039 : boolean := false;
    variable b1037 : boolean := false;
    variable b1035 : boolean := false;
    variable b1033 : boolean := false;
    variable b1031 : boolean := false;
    variable r1029 : std_logic_vector(0 to 31) := (others => '0');
    variable r1027 : std_logic_vector(0 to 31) := (others => '0');
    variable r1025 : std_logic_vector(0 to 31) := (others => '0');
    variable r1023 : std_logic_vector(0 to 31) := (others => '0');
    variable r1021 : std_logic_vector(0 to 31) := (others => '0');
    variable r1019 : std_logic_vector(0 to 31) := (others => '0');
    variable r1017 : std_logic_vector(0 to 31) := (others => '0');
    variable r1015 : std_logic_vector(0 to 31) := (others => '0');
    variable r1013 : std_logic_vector(0 to 31) := (others => '0');
    variable r1011 : std_logic_vector(0 to 31) := (others => '0');
    variable r1009 : std_logic_vector(0 to 31) := (others => '0');
    variable r1007 : std_logic_vector(0 to 31) := (others => '0');
    variable r1005 : std_logic_vector(0 to 31) := (others => '0');
    variable r1003 : std_logic_vector(0 to 31) := (others => '0');
    variable r1001 : std_logic_vector(0 to 31) := (others => '0');
    variable r999 : std_logic_vector(0 to 31) := (others => '0');
    variable b996 : boolean := false;
    variable b994 : boolean := false;
    variable r992 : std_logic_vector(0 to 511) := (others => '0');
    variable r990 : std_logic_vector(0 to 31) := (others => '0');
    variable r988 : std_logic_vector(0 to 31) := (others => '0');
    variable r986 : std_logic_vector(0 to 511) := (others => '0');
    variable r980 : std_logic_vector(0 to 575) := (others => '0');
    variable r977 : std_logic_vector(0 to 511) := (others => '0');
    variable b975 : boolean := false;
    variable b973 : boolean := false;
    variable b971 : boolean := false;
    variable r969 : std_logic_vector(0 to 31) := (others => '0');
    variable r967 : std_logic_vector(0 to 31) := (others => '0');
    variable b965 : boolean := false;
    variable r957 : std_logic_vector(0 to 67) := (others => '0');
    variable r953 : std_logic_vector(0 to 63) := (others => '0');
    variable r952 : std_logic_vector(0 to 64) := (others => '0');
    variable r950 : std_logic_vector(0 to 0) := (others => '0');
    variable r928 : std_logic_vector(0 to 511) := (others => '0');
    variable b925 : boolean := false;
    variable b923 : boolean := false;
    variable b921 : boolean := false;
    variable b919 : boolean := false;
    variable b917 : boolean := false;
    variable b915 : boolean := false;
    variable b913 : boolean := false;
    variable b911 : boolean := false;
    variable b909 : boolean := false;
    variable b907 : boolean := false;
    variable b905 : boolean := false;
    variable b903 : boolean := false;
    variable b901 : boolean := false;
    variable b899 : boolean := false;
    variable b897 : boolean := false;
    variable b895 : boolean := false;
    variable r893 : std_logic_vector(0 to 31) := (others => '0');
    variable r891 : std_logic_vector(0 to 31) := (others => '0');
    variable r889 : std_logic_vector(0 to 31) := (others => '0');
    variable r887 : std_logic_vector(0 to 31) := (others => '0');
    variable r885 : std_logic_vector(0 to 31) := (others => '0');
    variable r883 : std_logic_vector(0 to 31) := (others => '0');
    variable r881 : std_logic_vector(0 to 31) := (others => '0');
    variable r879 : std_logic_vector(0 to 31) := (others => '0');
    variable r877 : std_logic_vector(0 to 31) := (others => '0');
    variable r875 : std_logic_vector(0 to 31) := (others => '0');
    variable r873 : std_logic_vector(0 to 31) := (others => '0');
    variable r871 : std_logic_vector(0 to 31) := (others => '0');
    variable r869 : std_logic_vector(0 to 31) := (others => '0');
    variable r867 : std_logic_vector(0 to 31) := (others => '0');
    variable r865 : std_logic_vector(0 to 31) := (others => '0');
    variable r863 : std_logic_vector(0 to 31) := (others => '0');
    variable b860 : boolean := false;
    variable b858 : boolean := false;
    variable r856 : std_logic_vector(0 to 511) := (others => '0');
    variable r854 : std_logic_vector(0 to 31) := (others => '0');
    variable r852 : std_logic_vector(0 to 31) := (others => '0');
    variable r850 : std_logic_vector(0 to 511) := (others => '0');
    variable r844 : std_logic_vector(0 to 575) := (others => '0');
    variable r841 : std_logic_vector(0 to 511) := (others => '0');
    variable b839 : boolean := false;
    variable b837 : boolean := false;
    variable b835 : boolean := false;
    variable r833 : std_logic_vector(0 to 31) := (others => '0');
    variable r831 : std_logic_vector(0 to 31) := (others => '0');
    variable b829 : boolean := false;
    variable r821 : std_logic_vector(0 to 67) := (others => '0');
    variable r817 : std_logic_vector(0 to 63) := (others => '0');
    variable r816 : std_logic_vector(0 to 64) := (others => '0');
    variable r814 : std_logic_vector(0 to 0) := (others => '0');
    variable r792 : std_logic_vector(0 to 511) := (others => '0');
    variable b789 : boolean := false;
    variable b787 : boolean := false;
    variable b785 : boolean := false;
    variable b783 : boolean := false;
    variable b781 : boolean := false;
    variable b779 : boolean := false;
    variable b777 : boolean := false;
    variable b775 : boolean := false;
    variable b773 : boolean := false;
    variable b771 : boolean := false;
    variable b769 : boolean := false;
    variable b767 : boolean := false;
    variable b765 : boolean := false;
    variable b763 : boolean := false;
    variable b761 : boolean := false;
    variable b759 : boolean := false;
    variable r757 : std_logic_vector(0 to 31) := (others => '0');
    variable r755 : std_logic_vector(0 to 31) := (others => '0');
    variable r753 : std_logic_vector(0 to 31) := (others => '0');
    variable r751 : std_logic_vector(0 to 31) := (others => '0');
    variable r749 : std_logic_vector(0 to 31) := (others => '0');
    variable r747 : std_logic_vector(0 to 31) := (others => '0');
    variable r745 : std_logic_vector(0 to 31) := (others => '0');
    variable r743 : std_logic_vector(0 to 31) := (others => '0');
    variable r741 : std_logic_vector(0 to 31) := (others => '0');
    variable r739 : std_logic_vector(0 to 31) := (others => '0');
    variable r737 : std_logic_vector(0 to 31) := (others => '0');
    variable r735 : std_logic_vector(0 to 31) := (others => '0');
    variable r733 : std_logic_vector(0 to 31) := (others => '0');
    variable r731 : std_logic_vector(0 to 31) := (others => '0');
    variable r729 : std_logic_vector(0 to 31) := (others => '0');
    variable r727 : std_logic_vector(0 to 31) := (others => '0');
    variable b724 : boolean := false;
    variable b722 : boolean := false;
    variable r720 : std_logic_vector(0 to 511) := (others => '0');
    variable r718 : std_logic_vector(0 to 31) := (others => '0');
    variable r716 : std_logic_vector(0 to 31) := (others => '0');
    variable r714 : std_logic_vector(0 to 511) := (others => '0');
    variable r708 : std_logic_vector(0 to 575) := (others => '0');
    variable r705 : std_logic_vector(0 to 511) := (others => '0');
    variable b703 : boolean := false;
    variable b701 : boolean := false;
    variable b699 : boolean := false;
    variable r697 : std_logic_vector(0 to 31) := (others => '0');
    variable r695 : std_logic_vector(0 to 31) := (others => '0');
    variable b693 : boolean := false;
    variable r685 : std_logic_vector(0 to 67) := (others => '0');
    variable r681 : std_logic_vector(0 to 63) := (others => '0');
    variable r680 : std_logic_vector(0 to 64) := (others => '0');
    variable r678 : std_logic_vector(0 to 0) := (others => '0');
    variable r656 : std_logic_vector(0 to 511) := (others => '0');
    variable b653 : boolean := false;
    variable b651 : boolean := false;
    variable b649 : boolean := false;
    variable b647 : boolean := false;
    variable b645 : boolean := false;
    variable b643 : boolean := false;
    variable b641 : boolean := false;
    variable b639 : boolean := false;
    variable b637 : boolean := false;
    variable b635 : boolean := false;
    variable b633 : boolean := false;
    variable b631 : boolean := false;
    variable b629 : boolean := false;
    variable b627 : boolean := false;
    variable b625 : boolean := false;
    variable b623 : boolean := false;
    variable r621 : std_logic_vector(0 to 31) := (others => '0');
    variable r619 : std_logic_vector(0 to 31) := (others => '0');
    variable r617 : std_logic_vector(0 to 31) := (others => '0');
    variable r615 : std_logic_vector(0 to 31) := (others => '0');
    variable r613 : std_logic_vector(0 to 31) := (others => '0');
    variable r611 : std_logic_vector(0 to 31) := (others => '0');
    variable r609 : std_logic_vector(0 to 31) := (others => '0');
    variable r607 : std_logic_vector(0 to 31) := (others => '0');
    variable r605 : std_logic_vector(0 to 31) := (others => '0');
    variable r603 : std_logic_vector(0 to 31) := (others => '0');
    variable r601 : std_logic_vector(0 to 31) := (others => '0');
    variable r599 : std_logic_vector(0 to 31) := (others => '0');
    variable r597 : std_logic_vector(0 to 31) := (others => '0');
    variable r595 : std_logic_vector(0 to 31) := (others => '0');
    variable r593 : std_logic_vector(0 to 31) := (others => '0');
    variable r591 : std_logic_vector(0 to 31) := (others => '0');
    variable b588 : boolean := false;
    variable b586 : boolean := false;
    variable r584 : std_logic_vector(0 to 511) := (others => '0');
    variable r582 : std_logic_vector(0 to 31) := (others => '0');
    variable r580 : std_logic_vector(0 to 31) := (others => '0');
    variable r578 : std_logic_vector(0 to 511) := (others => '0');
    variable r572 : std_logic_vector(0 to 575) := (others => '0');
    variable r569 : std_logic_vector(0 to 511) := (others => '0');
    variable r566 : std_logic_vector(0 to 255) := (others => '0');
    variable b26 : boolean := false;
    variable b24 : boolean := false;
    variable b22 : boolean := false;
    variable r20 : std_logic_vector(0 to 31) := (others => '0');
    variable r18 : std_logic_vector(0 to 31) := (others => '0');
    variable b16 : boolean := false;
    variable r12 : std_logic_vector(0 to 67) := (others => '0');
    variable r10 : std_logic_vector(0 to 67) := (others => '0');
    variable r6 : std_logic_vector(0 to 63) := (others => '0');
    variable r5 : std_logic_vector(0 to 64) := (others => '0');
    variable r3 : std_logic_vector(0 to 0) := (others => '0');
    variable statevar0 : std_logic_vector(0 to 255) := (others => '0');
    variable statevar1 : std_logic_vector(0 to 511) := (others => '0');
    variable statevar2 : std_logic_vector(0 to 255) := (others => '0');
    variable statevar3 : std_logic_vector(0 to 5) := (others => '0');
    variable output_tmp : std_logic_vector(0 to 64);
  begin
    -- Read reg temps.
    control := control_flop;
    input_tmp := input_flop;
    goto_L7851 := goto_L7851_flop;
    goto_L7844 := goto_L7844_flop;
    goto_L7806 := goto_L7806_flop;
    goto_L7767 := goto_L7767_flop;
    goto_L7728 := goto_L7728_flop;
    goto_L7570 := goto_L7570_flop;
    goto_L7690 := goto_L7690_flop;
    goto_L7575 := goto_L7575_flop;
    goto_L1784 := goto_L1784_flop;
    goto_L1785 := goto_L1785_flop;
    goto_L1638 := goto_L1638_flop;
    goto_L1502 := goto_L1502_flop;
    goto_L1366 := goto_L1366_flop;
    goto_L1230 := goto_L1230_flop;
    goto_L1094 := goto_L1094_flop;
    goto_L958 := goto_L958_flop;
    goto_L822 := goto_L822_flop;
    goto_L686 := goto_L686_flop;
    goto_L11 := goto_L11_flop;
    goto_L13 := goto_L13_flop;
    goto_L690 := goto_L690_flop;
    goto_L826 := goto_L826_flop;
    goto_L962 := goto_L962_flop;
    goto_L1098 := goto_L1098_flop;
    goto_L1234 := goto_L1234_flop;
    goto_L1370 := goto_L1370_flop;
    goto_L1506 := goto_L1506_flop;
    goto_L1642 := goto_L1642_flop;
    goto_L7693 := goto_L7693_flop;
    goto_L7732 := goto_L7732_flop;
    goto_L7771 := goto_L7771_flop;
    goto_L7810 := goto_L7810_flop;
    goto_L7777 := goto_L7777_flop;
    goto_L7738 := goto_L7738_flop;
    goto_L7699 := goto_L7699_flop;
    goto_L1658 := goto_L1658_flop;
    goto_L1522 := goto_L1522_flop;
    goto_L1386 := goto_L1386_flop;
    goto_L1250 := goto_L1250_flop;
    goto_L1114 := goto_L1114_flop;
    goto_L978 := goto_L978_flop;
    goto_L842 := goto_L842_flop;
    goto_L706 := goto_L706_flop;
    goto_L567 := goto_L567_flop;
    goto_L0 := goto_L0_flop;
    goto_L7852 := goto_L7852_flop;
    r7843 := r7843_flop;
    r7840 := r7840_flop;
    r7817 := r7817_flop;
    r7814 := r7814_flop;
    r7805 := r7805_flop;
    r7802 := r7802_flop;
    r7779 := r7779_flop;
    r7776 := r7776_flop;
    b7774 := b7774_flop;
    r7766 := r7766_flop;
    r7763 := r7763_flop;
    r7740 := r7740_flop;
    r7737 := r7737_flop;
    b7735 := b7735_flop;
    r7727 := r7727_flop;
    r7724 := r7724_flop;
    r7701 := r7701_flop;
    r7698 := r7698_flop;
    b7696 := b7696_flop;
    r7679 := r7679_flop;
    r7675 := r7675_flop;
    r7671 := r7671_flop;
    r7667 := r7667_flop;
    r7663 := r7663_flop;
    r7659 := r7659_flop;
    r7655 := r7655_flop;
    r7651 := r7651_flop;
    r7647 := r7647_flop;
    b7644 := b7644_flop;
    b7642 := b7642_flop;
    b7640 := b7640_flop;
    b7638 := b7638_flop;
    b7636 := b7636_flop;
    b7634 := b7634_flop;
    b7632 := b7632_flop;
    b7630 := b7630_flop;
    r7628 := r7628_flop;
    r7626 := r7626_flop;
    r7624 := r7624_flop;
    r7622 := r7622_flop;
    r7620 := r7620_flop;
    r7618 := r7618_flop;
    r7616 := r7616_flop;
    r7614 := r7614_flop;
    r7610 := r7610_flop;
    b7608 := b7608_flop;
    b7606 := b7606_flop;
    b7604 := b7604_flop;
    b7602 := b7602_flop;
    b7600 := b7600_flop;
    b7598 := b7598_flop;
    b7596 := b7596_flop;
    b7594 := b7594_flop;
    r7592 := r7592_flop;
    r7590 := r7590_flop;
    r7588 := r7588_flop;
    r7586 := r7586_flop;
    r7584 := r7584_flop;
    r7582 := r7582_flop;
    r7580 := r7580_flop;
    r7578 := r7578_flop;
    r7574 := r7574_flop;
    b7572 := b7572_flop;
    r7569 := r7569_flop;
    r7565 := r7565_flop;
    r7564 := r7564_flop;
    r7562 := r7562_flop;
    r7558 := r7558_flop;
    r7300 := r7300_flop;
    r7296 := r7296_flop;
    r7292 := r7292_flop;
    r2874 := r2874_flop;
    r2376 := r2376_flop;
    r2375 := r2375_flop;
    r2374 := r2374_flop;
    r2371 := r2371_flop;
    r2365 := r2365_flop;
    r1862 := r1862_flop;
    b1859 := b1859_flop;
    b1857 := b1857_flop;
    b1855 := b1855_flop;
    b1853 := b1853_flop;
    b1851 := b1851_flop;
    b1849 := b1849_flop;
    b1847 := b1847_flop;
    b1845 := b1845_flop;
    b1843 := b1843_flop;
    b1841 := b1841_flop;
    b1839 := b1839_flop;
    b1837 := b1837_flop;
    b1835 := b1835_flop;
    b1833 := b1833_flop;
    b1831 := b1831_flop;
    b1829 := b1829_flop;
    r1827 := r1827_flop;
    r1825 := r1825_flop;
    r1823 := r1823_flop;
    r1821 := r1821_flop;
    r1819 := r1819_flop;
    r1817 := r1817_flop;
    r1815 := r1815_flop;
    r1813 := r1813_flop;
    r1811 := r1811_flop;
    r1809 := r1809_flop;
    r1807 := r1807_flop;
    r1805 := r1805_flop;
    r1803 := r1803_flop;
    r1801 := r1801_flop;
    r1799 := r1799_flop;
    r1797 := r1797_flop;
    r1795 := r1795_flop;
    r1792 := r1792_flop;
    r1790 := r1790_flop;
    r1787 := r1787_flop;
    r1783 := r1783_flop;
    r1779 := r1779_flop;
    r1778 := r1778_flop;
    r1776 := r1776_flop;
    r1754 := r1754_flop;
    b1751 := b1751_flop;
    b1749 := b1749_flop;
    b1747 := b1747_flop;
    b1745 := b1745_flop;
    b1743 := b1743_flop;
    b1741 := b1741_flop;
    b1739 := b1739_flop;
    b1737 := b1737_flop;
    b1735 := b1735_flop;
    b1733 := b1733_flop;
    b1731 := b1731_flop;
    b1729 := b1729_flop;
    b1727 := b1727_flop;
    b1725 := b1725_flop;
    b1723 := b1723_flop;
    b1721 := b1721_flop;
    r1719 := r1719_flop;
    r1717 := r1717_flop;
    r1715 := r1715_flop;
    r1713 := r1713_flop;
    r1711 := r1711_flop;
    r1709 := r1709_flop;
    r1707 := r1707_flop;
    r1705 := r1705_flop;
    r1703 := r1703_flop;
    r1701 := r1701_flop;
    r1699 := r1699_flop;
    r1697 := r1697_flop;
    r1695 := r1695_flop;
    r1693 := r1693_flop;
    r1691 := r1691_flop;
    r1689 := r1689_flop;
    b1686 := b1686_flop;
    b1684 := b1684_flop;
    r1682 := r1682_flop;
    r1680 := r1680_flop;
    r1678 := r1678_flop;
    r1676 := r1676_flop;
    r1670 := r1670_flop;
    r1667 := r1667_flop;
    r1663 := r1663_flop;
    r1659 := r1659_flop;
    r1657 := r1657_flop;
    b1655 := b1655_flop;
    b1653 := b1653_flop;
    b1651 := b1651_flop;
    r1649 := r1649_flop;
    r1647 := r1647_flop;
    b1645 := b1645_flop;
    r1637 := r1637_flop;
    r1633 := r1633_flop;
    r1632 := r1632_flop;
    r1630 := r1630_flop;
    r1608 := r1608_flop;
    b1605 := b1605_flop;
    b1603 := b1603_flop;
    b1601 := b1601_flop;
    b1599 := b1599_flop;
    b1597 := b1597_flop;
    b1595 := b1595_flop;
    b1593 := b1593_flop;
    b1591 := b1591_flop;
    b1589 := b1589_flop;
    b1587 := b1587_flop;
    b1585 := b1585_flop;
    b1583 := b1583_flop;
    b1581 := b1581_flop;
    b1579 := b1579_flop;
    b1577 := b1577_flop;
    b1575 := b1575_flop;
    r1573 := r1573_flop;
    r1571 := r1571_flop;
    r1569 := r1569_flop;
    r1567 := r1567_flop;
    r1565 := r1565_flop;
    r1563 := r1563_flop;
    r1561 := r1561_flop;
    r1559 := r1559_flop;
    r1557 := r1557_flop;
    r1555 := r1555_flop;
    r1553 := r1553_flop;
    r1551 := r1551_flop;
    r1549 := r1549_flop;
    r1547 := r1547_flop;
    r1545 := r1545_flop;
    r1543 := r1543_flop;
    b1540 := b1540_flop;
    b1538 := b1538_flop;
    r1536 := r1536_flop;
    r1534 := r1534_flop;
    r1532 := r1532_flop;
    r1530 := r1530_flop;
    r1524 := r1524_flop;
    r1521 := r1521_flop;
    b1519 := b1519_flop;
    b1517 := b1517_flop;
    b1515 := b1515_flop;
    r1513 := r1513_flop;
    r1511 := r1511_flop;
    b1509 := b1509_flop;
    r1501 := r1501_flop;
    r1497 := r1497_flop;
    r1496 := r1496_flop;
    r1494 := r1494_flop;
    r1472 := r1472_flop;
    b1469 := b1469_flop;
    b1467 := b1467_flop;
    b1465 := b1465_flop;
    b1463 := b1463_flop;
    b1461 := b1461_flop;
    b1459 := b1459_flop;
    b1457 := b1457_flop;
    b1455 := b1455_flop;
    b1453 := b1453_flop;
    b1451 := b1451_flop;
    b1449 := b1449_flop;
    b1447 := b1447_flop;
    b1445 := b1445_flop;
    b1443 := b1443_flop;
    b1441 := b1441_flop;
    b1439 := b1439_flop;
    r1437 := r1437_flop;
    r1435 := r1435_flop;
    r1433 := r1433_flop;
    r1431 := r1431_flop;
    r1429 := r1429_flop;
    r1427 := r1427_flop;
    r1425 := r1425_flop;
    r1423 := r1423_flop;
    r1421 := r1421_flop;
    r1419 := r1419_flop;
    r1417 := r1417_flop;
    r1415 := r1415_flop;
    r1413 := r1413_flop;
    r1411 := r1411_flop;
    r1409 := r1409_flop;
    r1407 := r1407_flop;
    b1404 := b1404_flop;
    b1402 := b1402_flop;
    r1400 := r1400_flop;
    r1398 := r1398_flop;
    r1396 := r1396_flop;
    r1394 := r1394_flop;
    r1388 := r1388_flop;
    r1385 := r1385_flop;
    b1383 := b1383_flop;
    b1381 := b1381_flop;
    b1379 := b1379_flop;
    r1377 := r1377_flop;
    r1375 := r1375_flop;
    b1373 := b1373_flop;
    r1365 := r1365_flop;
    r1361 := r1361_flop;
    r1360 := r1360_flop;
    r1358 := r1358_flop;
    r1336 := r1336_flop;
    b1333 := b1333_flop;
    b1331 := b1331_flop;
    b1329 := b1329_flop;
    b1327 := b1327_flop;
    b1325 := b1325_flop;
    b1323 := b1323_flop;
    b1321 := b1321_flop;
    b1319 := b1319_flop;
    b1317 := b1317_flop;
    b1315 := b1315_flop;
    b1313 := b1313_flop;
    b1311 := b1311_flop;
    b1309 := b1309_flop;
    b1307 := b1307_flop;
    b1305 := b1305_flop;
    b1303 := b1303_flop;
    r1301 := r1301_flop;
    r1299 := r1299_flop;
    r1297 := r1297_flop;
    r1295 := r1295_flop;
    r1293 := r1293_flop;
    r1291 := r1291_flop;
    r1289 := r1289_flop;
    r1287 := r1287_flop;
    r1285 := r1285_flop;
    r1283 := r1283_flop;
    r1281 := r1281_flop;
    r1279 := r1279_flop;
    r1277 := r1277_flop;
    r1275 := r1275_flop;
    r1273 := r1273_flop;
    r1271 := r1271_flop;
    b1268 := b1268_flop;
    b1266 := b1266_flop;
    r1264 := r1264_flop;
    r1262 := r1262_flop;
    r1260 := r1260_flop;
    r1258 := r1258_flop;
    r1252 := r1252_flop;
    r1249 := r1249_flop;
    b1247 := b1247_flop;
    b1245 := b1245_flop;
    b1243 := b1243_flop;
    r1241 := r1241_flop;
    r1239 := r1239_flop;
    b1237 := b1237_flop;
    r1229 := r1229_flop;
    r1225 := r1225_flop;
    r1224 := r1224_flop;
    r1222 := r1222_flop;
    r1200 := r1200_flop;
    b1197 := b1197_flop;
    b1195 := b1195_flop;
    b1193 := b1193_flop;
    b1191 := b1191_flop;
    b1189 := b1189_flop;
    b1187 := b1187_flop;
    b1185 := b1185_flop;
    b1183 := b1183_flop;
    b1181 := b1181_flop;
    b1179 := b1179_flop;
    b1177 := b1177_flop;
    b1175 := b1175_flop;
    b1173 := b1173_flop;
    b1171 := b1171_flop;
    b1169 := b1169_flop;
    b1167 := b1167_flop;
    r1165 := r1165_flop;
    r1163 := r1163_flop;
    r1161 := r1161_flop;
    r1159 := r1159_flop;
    r1157 := r1157_flop;
    r1155 := r1155_flop;
    r1153 := r1153_flop;
    r1151 := r1151_flop;
    r1149 := r1149_flop;
    r1147 := r1147_flop;
    r1145 := r1145_flop;
    r1143 := r1143_flop;
    r1141 := r1141_flop;
    r1139 := r1139_flop;
    r1137 := r1137_flop;
    r1135 := r1135_flop;
    b1132 := b1132_flop;
    b1130 := b1130_flop;
    r1128 := r1128_flop;
    r1126 := r1126_flop;
    r1124 := r1124_flop;
    r1122 := r1122_flop;
    r1116 := r1116_flop;
    r1113 := r1113_flop;
    b1111 := b1111_flop;
    b1109 := b1109_flop;
    b1107 := b1107_flop;
    r1105 := r1105_flop;
    r1103 := r1103_flop;
    b1101 := b1101_flop;
    r1093 := r1093_flop;
    r1089 := r1089_flop;
    r1088 := r1088_flop;
    r1086 := r1086_flop;
    r1064 := r1064_flop;
    b1061 := b1061_flop;
    b1059 := b1059_flop;
    b1057 := b1057_flop;
    b1055 := b1055_flop;
    b1053 := b1053_flop;
    b1051 := b1051_flop;
    b1049 := b1049_flop;
    b1047 := b1047_flop;
    b1045 := b1045_flop;
    b1043 := b1043_flop;
    b1041 := b1041_flop;
    b1039 := b1039_flop;
    b1037 := b1037_flop;
    b1035 := b1035_flop;
    b1033 := b1033_flop;
    b1031 := b1031_flop;
    r1029 := r1029_flop;
    r1027 := r1027_flop;
    r1025 := r1025_flop;
    r1023 := r1023_flop;
    r1021 := r1021_flop;
    r1019 := r1019_flop;
    r1017 := r1017_flop;
    r1015 := r1015_flop;
    r1013 := r1013_flop;
    r1011 := r1011_flop;
    r1009 := r1009_flop;
    r1007 := r1007_flop;
    r1005 := r1005_flop;
    r1003 := r1003_flop;
    r1001 := r1001_flop;
    r999 := r999_flop;
    b996 := b996_flop;
    b994 := b994_flop;
    r992 := r992_flop;
    r990 := r990_flop;
    r988 := r988_flop;
    r986 := r986_flop;
    r980 := r980_flop;
    r977 := r977_flop;
    b975 := b975_flop;
    b973 := b973_flop;
    b971 := b971_flop;
    r969 := r969_flop;
    r967 := r967_flop;
    b965 := b965_flop;
    r957 := r957_flop;
    r953 := r953_flop;
    r952 := r952_flop;
    r950 := r950_flop;
    r928 := r928_flop;
    b925 := b925_flop;
    b923 := b923_flop;
    b921 := b921_flop;
    b919 := b919_flop;
    b917 := b917_flop;
    b915 := b915_flop;
    b913 := b913_flop;
    b911 := b911_flop;
    b909 := b909_flop;
    b907 := b907_flop;
    b905 := b905_flop;
    b903 := b903_flop;
    b901 := b901_flop;
    b899 := b899_flop;
    b897 := b897_flop;
    b895 := b895_flop;
    r893 := r893_flop;
    r891 := r891_flop;
    r889 := r889_flop;
    r887 := r887_flop;
    r885 := r885_flop;
    r883 := r883_flop;
    r881 := r881_flop;
    r879 := r879_flop;
    r877 := r877_flop;
    r875 := r875_flop;
    r873 := r873_flop;
    r871 := r871_flop;
    r869 := r869_flop;
    r867 := r867_flop;
    r865 := r865_flop;
    r863 := r863_flop;
    b860 := b860_flop;
    b858 := b858_flop;
    r856 := r856_flop;
    r854 := r854_flop;
    r852 := r852_flop;
    r850 := r850_flop;
    r844 := r844_flop;
    r841 := r841_flop;
    b839 := b839_flop;
    b837 := b837_flop;
    b835 := b835_flop;
    r833 := r833_flop;
    r831 := r831_flop;
    b829 := b829_flop;
    r821 := r821_flop;
    r817 := r817_flop;
    r816 := r816_flop;
    r814 := r814_flop;
    r792 := r792_flop;
    b789 := b789_flop;
    b787 := b787_flop;
    b785 := b785_flop;
    b783 := b783_flop;
    b781 := b781_flop;
    b779 := b779_flop;
    b777 := b777_flop;
    b775 := b775_flop;
    b773 := b773_flop;
    b771 := b771_flop;
    b769 := b769_flop;
    b767 := b767_flop;
    b765 := b765_flop;
    b763 := b763_flop;
    b761 := b761_flop;
    b759 := b759_flop;
    r757 := r757_flop;
    r755 := r755_flop;
    r753 := r753_flop;
    r751 := r751_flop;
    r749 := r749_flop;
    r747 := r747_flop;
    r745 := r745_flop;
    r743 := r743_flop;
    r741 := r741_flop;
    r739 := r739_flop;
    r737 := r737_flop;
    r735 := r735_flop;
    r733 := r733_flop;
    r731 := r731_flop;
    r729 := r729_flop;
    r727 := r727_flop;
    b724 := b724_flop;
    b722 := b722_flop;
    r720 := r720_flop;
    r718 := r718_flop;
    r716 := r716_flop;
    r714 := r714_flop;
    r708 := r708_flop;
    r705 := r705_flop;
    b703 := b703_flop;
    b701 := b701_flop;
    b699 := b699_flop;
    r697 := r697_flop;
    r695 := r695_flop;
    b693 := b693_flop;
    r685 := r685_flop;
    r681 := r681_flop;
    r680 := r680_flop;
    r678 := r678_flop;
    r656 := r656_flop;
    b653 := b653_flop;
    b651 := b651_flop;
    b649 := b649_flop;
    b647 := b647_flop;
    b645 := b645_flop;
    b643 := b643_flop;
    b641 := b641_flop;
    b639 := b639_flop;
    b637 := b637_flop;
    b635 := b635_flop;
    b633 := b633_flop;
    b631 := b631_flop;
    b629 := b629_flop;
    b627 := b627_flop;
    b625 := b625_flop;
    b623 := b623_flop;
    r621 := r621_flop;
    r619 := r619_flop;
    r617 := r617_flop;
    r615 := r615_flop;
    r613 := r613_flop;
    r611 := r611_flop;
    r609 := r609_flop;
    r607 := r607_flop;
    r605 := r605_flop;
    r603 := r603_flop;
    r601 := r601_flop;
    r599 := r599_flop;
    r597 := r597_flop;
    r595 := r595_flop;
    r593 := r593_flop;
    r591 := r591_flop;
    b588 := b588_flop;
    b586 := b586_flop;
    r584 := r584_flop;
    r582 := r582_flop;
    r580 := r580_flop;
    r578 := r578_flop;
    r572 := r572_flop;
    r569 := r569_flop;
    r566 := r566_flop;
    b26 := b26_flop;
    b24 := b24_flop;
    b22 := b22_flop;
    r20 := r20_flop;
    r18 := r18_flop;
    b16 := b16_flop;
    r12 := r12_flop;
    r10 := r10_flop;
    r6 := r6_flop;
    r5 := r5_flop;
    r3 := r3_flop;
    statevar0 := statevar0_flop;
    statevar1 := statevar1_flop;
    statevar2 := statevar2_flop;
    statevar3 := statevar3_flop;
    output_tmp := (others => '0');
    -- Loop body.
    goto_L7851 := false;
    goto_L7844 := false;
    goto_L7806 := false;
    goto_L7767 := false;
    goto_L7728 := false;
    goto_L7570 := false;
    goto_L7690 := false;
    goto_L7575 := false;
    goto_L1784 := false;
    goto_L1785 := false;
    goto_L1638 := false;
    goto_L1502 := false;
    goto_L1366 := false;
    goto_L1230 := false;
    goto_L1094 := false;
    goto_L958 := false;
    goto_L822 := false;
    goto_L686 := false;
    goto_L11 := false;
    goto_L13 := false;
    goto_L690 := false;
    goto_L826 := false;
    goto_L962 := false;
    goto_L1098 := false;
    goto_L1234 := false;
    goto_L1370 := false;
    goto_L1506 := false;
    goto_L1642 := false;
    goto_L7693 := false;
    goto_L7732 := false;
    goto_L7771 := false;
    goto_L7810 := false;
    goto_L7777 := false;
    goto_L7738 := false;
    goto_L7699 := false;
    goto_L1658 := false;
    goto_L1522 := false;
    goto_L1386 := false;
    goto_L1250 := false;
    goto_L1114 := false;
    goto_L978 := false;
    goto_L842 := false;
    goto_L706 := false;
    goto_L567 := false;
    goto_L0 := false;
    goto_L7852 := false;
    null; -- label L7851
    -- ENTER
    goto_L0 := (control = STATE0);
    if (NOT goto_L0) then
      goto_L11 := (control = STATE11);
      if (NOT goto_L11) then
        goto_L686 := (control = STATE686);
        if (NOT goto_L686) then
          goto_L822 := (control = STATE822);
          if (NOT goto_L822) then
            goto_L958 := (control = STATE958);
            if (NOT goto_L958) then
              goto_L1094 := (control = STATE1094);
              if (NOT goto_L1094) then
                goto_L1230 := (control = STATE1230);
                if (NOT goto_L1230) then
                  goto_L1366 := (control = STATE1366);
                  if (NOT goto_L1366) then
                    goto_L1502 := (control = STATE1502);
                    if (NOT goto_L1502) then
                      goto_L1638 := (control = STATE1638);
                      if (NOT goto_L1638) then
                        goto_L1784 := (control = STATE1784);
                        if (NOT goto_L1784) then
                          goto_L7570 := (control = STATE7570);
                          if (NOT goto_L7570) then
                            goto_L7728 := (control = STATE7728);
                            if (NOT goto_L7728) then
                              goto_L7767 := (control = STATE7767);
                              if (NOT goto_L7767) then
                                goto_L7806 := (control = STATE7806);
                                if (NOT goto_L7806) then
                                  goto_L7844 := (control = STATE7844);
                                  null; -- label L7844
                                  r7843 := input_tmp;
                                  -- got i@26K in r7843
                                  r12 := r7843;
                                  goto_L13 := true;
                                end if;
                                goto_L13 := goto_L13;
                                if (NOT goto_L13) then
                                  null; -- label L7806
                                  r7805 := input_tmp;
                                  -- got i@26I in r7805
                                  r12 := r7805;
                                  goto_L13 := true;
                                end if;
                                goto_L13 := goto_L13;
                              end if;
                              goto_L13 := goto_L13;
                              if (NOT goto_L13) then
                                null; -- label L7767
                                r7766 := input_tmp;
                                -- got i@26G in r7766
                                r12 := r7766;
                                goto_L13 := true;
                              end if;
                              goto_L13 := goto_L13;
                            end if;
                            goto_L13 := goto_L13;
                            if (NOT goto_L13) then
                              null; -- label L7728
                              r7727 := input_tmp;
                              -- got i@26E in r7727
                              r12 := r7727;
                              goto_L13 := true;
                            end if;
                            goto_L13 := goto_L13;
                          end if;
                          goto_L13 := goto_L13;
                          if (NOT goto_L13) then
                            null; -- label L7570
                            r7569 := input_tmp;
                            -- got ctr@27C in r1787
                            b7572 := ("111111" = r1787(0 to 5));
                            goto_L7575 := b7572;
                            if (NOT goto_L7575) then
                              goto_L7690 := (NOT b7572);
                              null; -- label L7690
                              -- alt exit (no match)
                              goto_L1785 := true;
                            end if;
                            goto_L1785 := goto_L1785;
                            if (NOT goto_L1785) then
                              null; -- label L7575
                              r7574 := statevar2;
                              -- got $48@27E in r7574
                              -- final pat
                              r7578 := r7574(0 to 31);
                              r7580 := r7574(32 to 63);
                              r7582 := r7574(64 to 95);
                              r7584 := r7574(96 to 127);
                              r7586 := r7574(128 to 159);
                              r7588 := r7574(160 to 191);
                              r7590 := r7574(192 to 223);
                              r7592 := r7574(224 to 255);
                              b7594 := true;
                              b7596 := true;
                              b7598 := true;
                              b7600 := true;
                              b7602 := true;
                              b7604 := true;
                              b7606 := true;
                              b7608 := true;
                              r7610 := statevar0;
                              -- got $47@27N in r7610
                              -- final pat
                              r7614 := r7610(0 to 31);
                              r7616 := r7610(32 to 63);
                              r7618 := r7610(64 to 95);
                              r7620 := r7610(96 to 127);
                              r7622 := r7610(128 to 159);
                              r7624 := r7610(160 to 191);
                              r7626 := r7610(192 to 223);
                              r7628 := r7610(224 to 255);
                              b7630 := true;
                              b7632 := true;
                              b7634 := true;
                              b7636 := true;
                              b7638 := true;
                              b7640 := true;
                              b7642 := true;
                              b7644 := true;
                              null;
                              null;
                              -- got a@27O in r7614
                              -- got h1@27F in r7578
                              r7651 := w32Plus(r7614,r7578);
                              -- got b@27P in r7616
                              -- got h2@27G in r7580
                              r7655 := w32Plus(r7616,r7580);
                              -- got c@27Q in r7618
                              -- got h3@27H in r7582
                              r7659 := w32Plus(r7618,r7582);
                              -- got d@27R in r7620
                              -- got h4@27I in r7584
                              r7663 := w32Plus(r7620,r7584);
                              -- got e@27S in r7622
                              -- got h5@27J in r7586
                              r7667 := w32Plus(r7622,r7586);
                              -- got f@27T in r7624
                              -- got h6@27K in r7588
                              r7671 := w32Plus(r7624,r7588);
                              -- got g@27U in r7626
                              -- got h7@27L in r7590
                              r7675 := w32Plus(r7626,r7590);
                              -- got h@27V in r7628
                              -- got h8@27M in r7592
                              r7679 := w32Plus(r7628,r7592);
                              r7647 := (r7651 & r7655 & r7659 & r7663 & r7667 & r7671 & r7675 & r7679);
                              statevar2 := r7647;
                              null;
                              -- end case
                              null;
                              -- end case
                              -- got i@27D in r7569
                              r12 := r7569;
                              goto_L13 := true;
                            end if;
                            goto_L13 := goto_L13;
                          end if;
                          goto_L13 := goto_L13;
                          if (NOT goto_L13) then
                            goto_L1785 := goto_L1785;
                          end if;
                          goto_L1785 := goto_L1785;
                        end if;
                        goto_L1785 := goto_L1785;
                        if (NOT goto_L1785) then
                          goto_L13 := goto_L13;
                          if (NOT goto_L13) then
                            null; -- label L1784
                            r1783 := input_tmp;
                            goto_L1785 := true;
                          end if;
                          goto_L1785 := goto_L1785;
                        end if;
                        goto_L1785 := goto_L1785;
                        if (NOT goto_L1785) then
                          goto_L13 := goto_L13;
                        end if;
                        goto_L13 := goto_L13;
                        if (NOT goto_L13) then
                          null; -- label L1785
                          -- Mainloop in
                          -- Maingenhash' in
                          r1790 := statevar3;
                          r1792 := statevar1;
                          -- got s@26M in r1792
                          -- final pat
                          r1797 := r1792(0 to 31);
                          r1799 := r1792(32 to 63);
                          r1801 := r1792(64 to 95);
                          r1803 := r1792(96 to 127);
                          r1805 := r1792(128 to 159);
                          r1807 := r1792(160 to 191);
                          r1809 := r1792(192 to 223);
                          r1811 := r1792(224 to 255);
                          r1813 := r1792(256 to 287);
                          r1815 := r1792(288 to 319);
                          r1817 := r1792(320 to 351);
                          r1819 := r1792(352 to 383);
                          r1821 := r1792(384 to 415);
                          r1823 := r1792(416 to 447);
                          r1825 := r1792(448 to 479);
                          r1827 := r1792(480 to 511);
                          b1829 := true;
                          b1831 := true;
                          b1833 := true;
                          b1835 := true;
                          b1837 := true;
                          b1839 := true;
                          b1841 := true;
                          b1843 := true;
                          b1845 := true;
                          b1847 := true;
                          b1849 := true;
                          b1851 := true;
                          b1853 := true;
                          b1855 := true;
                          b1857 := true;
                          b1859 := true;
                          -- got s@26M in r1792
                          r2365 := rewire_MainupdateSched_1861(r1792);
                          statevar1 := r2365;
                          -- got w00@26N in r1797
                          r1795 := r1797;
                          -- end case
                          r2371 := statevar0;
                          -- got ctr@26L in r1790
                          r7292 := rewire_Mainseed_2873(r1790);
                          -- got $12@278 in r1795
                          -- got s@279 in r2371
                          r7296 := rewire_Mainstep256_2373(r7292,r1795,r2371);
                          statevar0 := r7296;
                          -- got ctr@26L in r1790
                          r7558 := rewire_MainincCtr_7299(r1790);
                          statevar3 := r7558;
                          -- got ctr@26L in r1790
                          -- Maingenhash' out
                          r7562 := "1";
                          r7565 := "0000000000000000000000000000000000000000000000000000000000000000";
                          r7564 := (r7562 & r7565);
                          output_tmp := r7564;
                          control := STATE7570;
                          goto_L7852 := true;
                        end if;
                        goto_L7852 := goto_L7852;
                      end if;
                      goto_L7852 := goto_L7852;
                      if (NOT goto_L7852) then
                        goto_L13 := goto_L13;
                        if (NOT goto_L13) then
                          null; -- label L1638
                          r1637 := input_tmp;
                          -- got i@25I in r1637
                          r12 := r1637;
                          goto_L13 := true;
                        end if;
                        goto_L13 := goto_L13;
                      end if;
                      goto_L13 := goto_L13;
                    end if;
                    goto_L13 := goto_L13;
                    if (NOT goto_L13) then
                      goto_L7852 := goto_L7852;
                      if (NOT goto_L7852) then
                        null; -- label L1502
                        r1501 := input_tmp;
                        -- got i@24R in r1501
                        r12 := r1501;
                        goto_L13 := true;
                      end if;
                      goto_L13 := goto_L13;
                    end if;
                    goto_L13 := goto_L13;
                    if (NOT goto_L13) then
                      goto_L7852 := goto_L7852;
                    end if;
                    goto_L7852 := goto_L7852;
                  end if;
                  goto_L7852 := goto_L7852;
                  if (NOT goto_L7852) then
                    goto_L13 := goto_L13;
                    if (NOT goto_L13) then
                      null; -- label L1366
                      r1365 := input_tmp;
                      -- got i@244 in r1365
                      r12 := r1365;
                      goto_L13 := true;
                    end if;
                    goto_L13 := goto_L13;
                  end if;
                  goto_L13 := goto_L13;
                end if;
                goto_L13 := goto_L13;
                if (NOT goto_L13) then
                  goto_L7852 := goto_L7852;
                  if (NOT goto_L7852) then
                    null; -- label L1230
                    r1229 := input_tmp;
                    -- got i@23D in r1229
                    r12 := r1229;
                    goto_L13 := true;
                  end if;
                  goto_L13 := goto_L13;
                end if;
                goto_L13 := goto_L13;
                if (NOT goto_L13) then
                  goto_L7852 := goto_L7852;
                end if;
                goto_L7852 := goto_L7852;
              end if;
              goto_L7852 := goto_L7852;
              if (NOT goto_L7852) then
                goto_L13 := goto_L13;
                if (NOT goto_L13) then
                  null; -- label L1094
                  r1093 := input_tmp;
                  -- got i@22M in r1093
                  r12 := r1093;
                  goto_L13 := true;
                end if;
                goto_L13 := goto_L13;
              end if;
              goto_L13 := goto_L13;
            end if;
            goto_L13 := goto_L13;
            if (NOT goto_L13) then
              goto_L7852 := goto_L7852;
              if (NOT goto_L7852) then
                null; -- label L958
                r957 := input_tmp;
                -- got i@21V in r957
                r12 := r957;
                goto_L13 := true;
              end if;
              goto_L13 := goto_L13;
            end if;
            goto_L13 := goto_L13;
            if (NOT goto_L13) then
              goto_L7852 := goto_L7852;
            end if;
            goto_L7852 := goto_L7852;
          end if;
          goto_L7852 := goto_L7852;
          if (NOT goto_L7852) then
            goto_L13 := goto_L13;
            if (NOT goto_L13) then
              null; -- label L822
              r821 := input_tmp;
              -- got i@218 in r821
              r12 := r821;
              goto_L13 := true;
            end if;
            goto_L13 := goto_L13;
          end if;
          goto_L13 := goto_L13;
        end if;
        goto_L13 := goto_L13;
        if (NOT goto_L13) then
          goto_L7852 := goto_L7852;
          if (NOT goto_L7852) then
            null; -- label L686
            r685 := input_tmp;
            -- got i@20H in r685
            r12 := r685;
            goto_L13 := true;
          end if;
          goto_L13 := goto_L13;
        end if;
        goto_L13 := goto_L13;
        if (NOT goto_L13) then
          goto_L7852 := goto_L7852;
        end if;
        goto_L7852 := goto_L7852;
      end if;
      goto_L7852 := goto_L7852;
      if (NOT goto_L7852) then
        goto_L13 := goto_L13;
        if (NOT goto_L13) then
          null; -- label L11
          r10 := input_tmp;
          -- got d@1VO in r10
          r12 := r10;
          goto_L13 := true;
        end if;
        goto_L13 := goto_L13;
        null; -- label L13
        -- Maindev in
        -- got $44@1VP in r12
        b16 := ("0000" = r12(0 to 3));
        r18 := r12(4 to 35);
        r20 := r12(36 to 67);
        b22 := true;
        b24 := true;
        b26 := (b16 AND (b22 AND b24));
        goto_L567 := b26;
        if (NOT goto_L567) then
          goto_L690 := (NOT b26);
          null; -- label L690
          -- alt exit (no match)
          -- got $44@1VP in r12
          b693 := ("0001" = r12(0 to 3));
          r695 := r12(4 to 35);
          r697 := r12(36 to 67);
          b699 := true;
          b701 := true;
          b703 := (b693 AND (b699 AND b701));
          goto_L706 := b703;
          if (NOT goto_L706) then
            goto_L826 := (NOT b703);
            null; -- label L826
            -- alt exit (no match)
            -- got $44@1VP in r12
            b829 := ("0010" = r12(0 to 3));
            r831 := r12(4 to 35);
            r833 := r12(36 to 67);
            b835 := true;
            b837 := true;
            b839 := (b829 AND (b835 AND b837));
            goto_L842 := b839;
            if (NOT goto_L842) then
              goto_L962 := (NOT b839);
              null; -- label L962
              -- alt exit (no match)
              -- got $44@1VP in r12
              b965 := ("0011" = r12(0 to 3));
              r967 := r12(4 to 35);
              r969 := r12(36 to 67);
              b971 := true;
              b973 := true;
              b975 := (b965 AND (b971 AND b973));
              goto_L978 := b975;
              if (NOT goto_L978) then
                goto_L1098 := (NOT b975);
                null; -- label L1098
                -- alt exit (no match)
                -- got $44@1VP in r12
                b1101 := ("0100" = r12(0 to 3));
                r1103 := r12(4 to 35);
                r1105 := r12(36 to 67);
                b1107 := true;
                b1109 := true;
                b1111 := (b1101 AND (b1107 AND b1109));
                goto_L1114 := b1111;
                if (NOT goto_L1114) then
                  goto_L1234 := (NOT b1111);
                  null; -- label L1234
                  -- alt exit (no match)
                  -- got $44@1VP in r12
                  b1237 := ("0101" = r12(0 to 3));
                  r1239 := r12(4 to 35);
                  r1241 := r12(36 to 67);
                  b1243 := true;
                  b1245 := true;
                  b1247 := (b1237 AND (b1243 AND b1245));
                  goto_L1250 := b1247;
                  if (NOT goto_L1250) then
                    goto_L1370 := (NOT b1247);
                    null; -- label L1370
                    -- alt exit (no match)
                    -- got $44@1VP in r12
                    b1373 := ("0110" = r12(0 to 3));
                    r1375 := r12(4 to 35);
                    r1377 := r12(36 to 67);
                    b1379 := true;
                    b1381 := true;
                    b1383 := (b1373 AND (b1379 AND b1381));
                    goto_L1386 := b1383;
                    if (NOT goto_L1386) then
                      goto_L1506 := (NOT b1383);
                      null; -- label L1506
                      -- alt exit (no match)
                      -- got $44@1VP in r12
                      b1509 := ("0111" = r12(0 to 3));
                      r1511 := r12(4 to 35);
                      r1513 := r12(36 to 67);
                      b1515 := true;
                      b1517 := true;
                      b1519 := (b1509 AND (b1515 AND b1517));
                      goto_L1522 := b1519;
                      if (NOT goto_L1522) then
                        goto_L1642 := (NOT b1519);
                        null; -- label L1642
                        -- alt exit (no match)
                        -- got $44@1VP in r12
                        b1645 := ("1000" = r12(0 to 3));
                        r1647 := r12(4 to 35);
                        r1649 := r12(36 to 67);
                        b1651 := true;
                        b1653 := true;
                        b1655 := (b1645 AND (b1651 AND b1653));
                        goto_L1658 := b1655;
                        if (NOT goto_L1658) then
                          goto_L7693 := (NOT b1655);
                          null; -- label L7693
                          -- alt exit (no match)
                          -- got $44@1VP in r12
                          b7696 := ("1001" = r12(0 to 3));
                          goto_L7699 := b7696;
                          if (NOT goto_L7699) then
                            goto_L7732 := (NOT b7696);
                            null; -- label L7732
                            -- alt exit (no match)
                            -- got $44@1VP in r12
                            b7735 := ("1010" = r12(0 to 3));
                            goto_L7738 := b7735;
                            if (NOT goto_L7738) then
                              goto_L7771 := (NOT b7735);
                              null; -- label L7771
                              -- alt exit (no match)
                              -- got $44@1VP in r12
                              b7774 := ("1011" = r12(0 to 3));
                              goto_L7777 := b7774;
                              if (NOT goto_L7777) then
                                goto_L7810 := (NOT b7774);
                                null; -- label L7810
                                -- alt exit (no match)
                                -- got $44@1VP in r12
                                -- final pat
                                r7814 := statevar2;
                                -- got h_n@26J in r7814
                                r7840 := rewire_Maindigest3_7816(r7814);
                                output_tmp := r7840;
                                control := STATE7844;
                                goto_L7852 := true;
                              end if;
                              goto_L7852 := goto_L7852;
                              if (NOT goto_L7852) then
                                null; -- label L7777
                                r7776 := statevar2;
                                -- got h_n@26H in r7776
                                r7802 := rewire_Maindigest2_7778(r7776);
                                output_tmp := r7802;
                                control := STATE7806;
                                goto_L7852 := true;
                              end if;
                              goto_L7852 := goto_L7852;
                            end if;
                            goto_L7852 := goto_L7852;
                            if (NOT goto_L7852) then
                              null; -- label L7738
                              r7737 := statevar2;
                              -- got h_n@26F in r7737
                              r7763 := rewire_Maindigest1_7739(r7737);
                              output_tmp := r7763;
                              control := STATE7767;
                              goto_L7852 := true;
                            end if;
                            goto_L7852 := goto_L7852;
                          end if;
                          goto_L7852 := goto_L7852;
                          if (NOT goto_L7852) then
                            null; -- label L7699
                            r7698 := statevar2;
                            -- got h_n@26D in r7698
                            r7724 := rewire_Maindigest0_7700(r7698);
                            output_tmp := r7724;
                            control := STATE7728;
                            goto_L7852 := true;
                          end if;
                          goto_L7852 := goto_L7852;
                        end if;
                        goto_L7852 := goto_L7852;
                        if (NOT goto_L7852) then
                          null; -- label L1658
                          r1657 := "000000";
                          null;
                          r1659 := (r1657);
                          statevar3 := r1659;
                          r1663 := statevar2;
                          -- got hi_1@25M in r1663
                          statevar0 := r1663;
                          r1667 := statevar1;
                          null;
                          null;
                          -- got w1@25J in r1647
                          -- got w2@25K in r1649
                          -- got hw@25O in r1667
                          r1670 := (r1647 & r1649 & r1667);
                          -- final pat
                          r1678 := r1670(0 to 31);
                          r1680 := r1670(32 to 63);
                          r1682 := r1670(64 to 575);
                          b1684 := true;
                          b1686 := true;
                          -- final pat
                          r1689 := r1682(0 to 31);
                          r1691 := r1682(32 to 63);
                          r1693 := r1682(64 to 95);
                          r1695 := r1682(96 to 127);
                          r1697 := r1682(128 to 159);
                          r1699 := r1682(160 to 191);
                          r1701 := r1682(192 to 223);
                          r1703 := r1682(224 to 255);
                          r1705 := r1682(256 to 287);
                          r1707 := r1682(288 to 319);
                          r1709 := r1682(320 to 351);
                          r1711 := r1682(352 to 383);
                          r1713 := r1682(384 to 415);
                          r1715 := r1682(416 to 447);
                          r1717 := r1682(448 to 479);
                          r1719 := r1682(480 to 511);
                          b1721 := true;
                          b1723 := true;
                          b1725 := true;
                          b1727 := true;
                          b1729 := true;
                          b1731 := true;
                          b1733 := true;
                          b1735 := true;
                          b1737 := true;
                          b1739 := true;
                          b1741 := true;
                          b1743 := true;
                          b1745 := true;
                          b1747 := true;
                          b1749 := true;
                          b1751 := true;
                          null;
                          null;
                          -- got x0@25R in r1689
                          -- got x1@25S in r1691
                          -- got x2@25T in r1693
                          -- got x3@25U in r1695
                          -- got x4@25V in r1697
                          -- got x5@260 in r1699
                          -- got x6@261 in r1701
                          -- got x7@262 in r1703
                          -- got x8@263 in r1705
                          -- got x9@264 in r1707
                          -- got xa@265 in r1709
                          -- got xb@266 in r1711
                          -- got xc@267 in r1713
                          -- got xd@268 in r1715
                          -- got w1'@25P in r1678
                          -- got w2'@25Q in r1680
                          r1754 := (r1689 & r1691 & r1693 & r1695 & r1697 & r1699 & r1701 & r1703 & r1705 & r1707 & r1709 & r1711 & r1713 & r1715 & r1678 & r1680);
                          r1676 := r1754;
                          -- end case
                          statevar1 := r1676;
                          r1776 := "1";
                          r1779 := "0000000000000000000000000000000000000000000000000000000000000000";
                          r1778 := (r1776 & r1779);
                          output_tmp := r1778;
                          control := STATE1784;
                          goto_L7852 := true;
                        end if;
                        goto_L7852 := goto_L7852;
                      end if;
                      goto_L7852 := goto_L7852;
                      if (NOT goto_L7852) then
                        null; -- label L1522
                        r1521 := statevar1;
                        null;
                        null;
                        -- got w1@24S in r1511
                        -- got w2@24T in r1513
                        -- got hw@24U in r1521
                        r1524 := (r1511 & r1513 & r1521);
                        -- final pat
                        r1532 := r1524(0 to 31);
                        r1534 := r1524(32 to 63);
                        r1536 := r1524(64 to 575);
                        b1538 := true;
                        b1540 := true;
                        -- final pat
                        r1543 := r1536(0 to 31);
                        r1545 := r1536(32 to 63);
                        r1547 := r1536(64 to 95);
                        r1549 := r1536(96 to 127);
                        r1551 := r1536(128 to 159);
                        r1553 := r1536(160 to 191);
                        r1555 := r1536(192 to 223);
                        r1557 := r1536(224 to 255);
                        r1559 := r1536(256 to 287);
                        r1561 := r1536(288 to 319);
                        r1563 := r1536(320 to 351);
                        r1565 := r1536(352 to 383);
                        r1567 := r1536(384 to 415);
                        r1569 := r1536(416 to 447);
                        r1571 := r1536(448 to 479);
                        r1573 := r1536(480 to 511);
                        b1575 := true;
                        b1577 := true;
                        b1579 := true;
                        b1581 := true;
                        b1583 := true;
                        b1585 := true;
                        b1587 := true;
                        b1589 := true;
                        b1591 := true;
                        b1593 := true;
                        b1595 := true;
                        b1597 := true;
                        b1599 := true;
                        b1601 := true;
                        b1603 := true;
                        b1605 := true;
                        null;
                        null;
                        -- got x0@251 in r1543
                        -- got x1@252 in r1545
                        -- got x2@253 in r1547
                        -- got x3@254 in r1549
                        -- got x4@255 in r1551
                        -- got x5@256 in r1553
                        -- got x6@257 in r1555
                        -- got x7@258 in r1557
                        -- got x8@259 in r1559
                        -- got x9@25A in r1561
                        -- got xa@25B in r1563
                        -- got xb@25C in r1565
                        -- got w1'@24V in r1532
                        -- got w2'@250 in r1534
                        -- got xe@25F in r1571
                        -- got xf@25G in r1573
                        r1608 := (r1543 & r1545 & r1547 & r1549 & r1551 & r1553 & r1555 & r1557 & r1559 & r1561 & r1563 & r1565 & r1532 & r1534 & r1571 & r1573);
                        r1530 := r1608;
                        -- end case
                        statevar1 := r1530;
                        r1630 := "1";
                        r1633 := "0000000000000000000000000000000000000000000000000000000000000000";
                        r1632 := (r1630 & r1633);
                        output_tmp := r1632;
                        control := STATE1638;
                        goto_L7852 := true;
                      end if;
                      goto_L7852 := goto_L7852;
                    end if;
                    goto_L7852 := goto_L7852;
                    if (NOT goto_L7852) then
                      null; -- label L1386
                      r1385 := statevar1;
                      null;
                      null;
                      -- got w1@245 in r1375
                      -- got w2@246 in r1377
                      -- got hw@247 in r1385
                      r1388 := (r1375 & r1377 & r1385);
                      -- final pat
                      r1396 := r1388(0 to 31);
                      r1398 := r1388(32 to 63);
                      r1400 := r1388(64 to 575);
                      b1402 := true;
                      b1404 := true;
                      -- final pat
                      r1407 := r1400(0 to 31);
                      r1409 := r1400(32 to 63);
                      r1411 := r1400(64 to 95);
                      r1413 := r1400(96 to 127);
                      r1415 := r1400(128 to 159);
                      r1417 := r1400(160 to 191);
                      r1419 := r1400(192 to 223);
                      r1421 := r1400(224 to 255);
                      r1423 := r1400(256 to 287);
                      r1425 := r1400(288 to 319);
                      r1427 := r1400(320 to 351);
                      r1429 := r1400(352 to 383);
                      r1431 := r1400(384 to 415);
                      r1433 := r1400(416 to 447);
                      r1435 := r1400(448 to 479);
                      r1437 := r1400(480 to 511);
                      b1439 := true;
                      b1441 := true;
                      b1443 := true;
                      b1445 := true;
                      b1447 := true;
                      b1449 := true;
                      b1451 := true;
                      b1453 := true;
                      b1455 := true;
                      b1457 := true;
                      b1459 := true;
                      b1461 := true;
                      b1463 := true;
                      b1465 := true;
                      b1467 := true;
                      b1469 := true;
                      null;
                      null;
                      -- got x0@24A in r1407
                      -- got x1@24B in r1409
                      -- got x2@24C in r1411
                      -- got x3@24D in r1413
                      -- got x4@24E in r1415
                      -- got x5@24F in r1417
                      -- got x6@24G in r1419
                      -- got x7@24H in r1421
                      -- got x8@24I in r1423
                      -- got x9@24J in r1425
                      -- got w1'@248 in r1396
                      -- got w2'@249 in r1398
                      -- got xc@24M in r1431
                      -- got xd@24N in r1433
                      -- got xe@24O in r1435
                      -- got xf@24P in r1437
                      r1472 := (r1407 & r1409 & r1411 & r1413 & r1415 & r1417 & r1419 & r1421 & r1423 & r1425 & r1396 & r1398 & r1431 & r1433 & r1435 & r1437);
                      r1394 := r1472;
                      -- end case
                      statevar1 := r1394;
                      r1494 := "1";
                      r1497 := "0000000000000000000000000000000000000000000000000000000000000000";
                      r1496 := (r1494 & r1497);
                      output_tmp := r1496;
                      control := STATE1502;
                      goto_L7852 := true;
                    end if;
                    goto_L7852 := goto_L7852;
                  end if;
                  goto_L7852 := goto_L7852;
                  if (NOT goto_L7852) then
                    null; -- label L1250
                    r1249 := statevar1;
                    null;
                    null;
                    -- got w1@23E in r1239
                    -- got w2@23F in r1241
                    -- got hw@23G in r1249
                    r1252 := (r1239 & r1241 & r1249);
                    -- final pat
                    r1260 := r1252(0 to 31);
                    r1262 := r1252(32 to 63);
                    r1264 := r1252(64 to 575);
                    b1266 := true;
                    b1268 := true;
                    -- final pat
                    r1271 := r1264(0 to 31);
                    r1273 := r1264(32 to 63);
                    r1275 := r1264(64 to 95);
                    r1277 := r1264(96 to 127);
                    r1279 := r1264(128 to 159);
                    r1281 := r1264(160 to 191);
                    r1283 := r1264(192 to 223);
                    r1285 := r1264(224 to 255);
                    r1287 := r1264(256 to 287);
                    r1289 := r1264(288 to 319);
                    r1291 := r1264(320 to 351);
                    r1293 := r1264(352 to 383);
                    r1295 := r1264(384 to 415);
                    r1297 := r1264(416 to 447);
                    r1299 := r1264(448 to 479);
                    r1301 := r1264(480 to 511);
                    b1303 := true;
                    b1305 := true;
                    b1307 := true;
                    b1309 := true;
                    b1311 := true;
                    b1313 := true;
                    b1315 := true;
                    b1317 := true;
                    b1319 := true;
                    b1321 := true;
                    b1323 := true;
                    b1325 := true;
                    b1327 := true;
                    b1329 := true;
                    b1331 := true;
                    b1333 := true;
                    null;
                    null;
                    -- got x0@23J in r1271
                    -- got x1@23K in r1273
                    -- got x2@23L in r1275
                    -- got x3@23M in r1277
                    -- got x4@23N in r1279
                    -- got x5@23O in r1281
                    -- got x6@23P in r1283
                    -- got x7@23Q in r1285
                    -- got w1'@23H in r1260
                    -- got w2'@23I in r1262
                    -- got xa@23T in r1291
                    -- got xb@23U in r1293
                    -- got xc@23V in r1295
                    -- got xd@240 in r1297
                    -- got xe@241 in r1299
                    -- got xf@242 in r1301
                    r1336 := (r1271 & r1273 & r1275 & r1277 & r1279 & r1281 & r1283 & r1285 & r1260 & r1262 & r1291 & r1293 & r1295 & r1297 & r1299 & r1301);
                    r1258 := r1336;
                    -- end case
                    statevar1 := r1258;
                    r1358 := "1";
                    r1361 := "0000000000000000000000000000000000000000000000000000000000000000";
                    r1360 := (r1358 & r1361);
                    output_tmp := r1360;
                    control := STATE1366;
                    goto_L7852 := true;
                  end if;
                  goto_L7852 := goto_L7852;
                end if;
                goto_L7852 := goto_L7852;
                if (NOT goto_L7852) then
                  null; -- label L1114
                  r1113 := statevar1;
                  null;
                  null;
                  -- got w1@22N in r1103
                  -- got w2@22O in r1105
                  -- got hw@22P in r1113
                  r1116 := (r1103 & r1105 & r1113);
                  -- final pat
                  r1124 := r1116(0 to 31);
                  r1126 := r1116(32 to 63);
                  r1128 := r1116(64 to 575);
                  b1130 := true;
                  b1132 := true;
                  -- final pat
                  r1135 := r1128(0 to 31);
                  r1137 := r1128(32 to 63);
                  r1139 := r1128(64 to 95);
                  r1141 := r1128(96 to 127);
                  r1143 := r1128(128 to 159);
                  r1145 := r1128(160 to 191);
                  r1147 := r1128(192 to 223);
                  r1149 := r1128(224 to 255);
                  r1151 := r1128(256 to 287);
                  r1153 := r1128(288 to 319);
                  r1155 := r1128(320 to 351);
                  r1157 := r1128(352 to 383);
                  r1159 := r1128(384 to 415);
                  r1161 := r1128(416 to 447);
                  r1163 := r1128(448 to 479);
                  r1165 := r1128(480 to 511);
                  b1167 := true;
                  b1169 := true;
                  b1171 := true;
                  b1173 := true;
                  b1175 := true;
                  b1177 := true;
                  b1179 := true;
                  b1181 := true;
                  b1183 := true;
                  b1185 := true;
                  b1187 := true;
                  b1189 := true;
                  b1191 := true;
                  b1193 := true;
                  b1195 := true;
                  b1197 := true;
                  null;
                  null;
                  -- got x0@22S in r1135
                  -- got x1@22T in r1137
                  -- got x2@22U in r1139
                  -- got x3@22V in r1141
                  -- got x4@230 in r1143
                  -- got x5@231 in r1145
                  -- got w1'@22Q in r1124
                  -- got w2'@22R in r1126
                  -- got x8@234 in r1151
                  -- got x9@235 in r1153
                  -- got xa@236 in r1155
                  -- got xb@237 in r1157
                  -- got xc@238 in r1159
                  -- got xd@239 in r1161
                  -- got xe@23A in r1163
                  -- got xf@23B in r1165
                  r1200 := (r1135 & r1137 & r1139 & r1141 & r1143 & r1145 & r1124 & r1126 & r1151 & r1153 & r1155 & r1157 & r1159 & r1161 & r1163 & r1165);
                  r1122 := r1200;
                  -- end case
                  statevar1 := r1122;
                  r1222 := "1";
                  r1225 := "0000000000000000000000000000000000000000000000000000000000000000";
                  r1224 := (r1222 & r1225);
                  output_tmp := r1224;
                  control := STATE1230;
                  goto_L7852 := true;
                end if;
                goto_L7852 := goto_L7852;
              end if;
              goto_L7852 := goto_L7852;
              if (NOT goto_L7852) then
                null; -- label L978
                r977 := statevar1;
                null;
                null;
                -- got w1@220 in r967
                -- got w2@221 in r969
                -- got hw@222 in r977
                r980 := (r967 & r969 & r977);
                -- final pat
                r988 := r980(0 to 31);
                r990 := r980(32 to 63);
                r992 := r980(64 to 575);
                b994 := true;
                b996 := true;
                -- final pat
                r999 := r992(0 to 31);
                r1001 := r992(32 to 63);
                r1003 := r992(64 to 95);
                r1005 := r992(96 to 127);
                r1007 := r992(128 to 159);
                r1009 := r992(160 to 191);
                r1011 := r992(192 to 223);
                r1013 := r992(224 to 255);
                r1015 := r992(256 to 287);
                r1017 := r992(288 to 319);
                r1019 := r992(320 to 351);
                r1021 := r992(352 to 383);
                r1023 := r992(384 to 415);
                r1025 := r992(416 to 447);
                r1027 := r992(448 to 479);
                r1029 := r992(480 to 511);
                b1031 := true;
                b1033 := true;
                b1035 := true;
                b1037 := true;
                b1039 := true;
                b1041 := true;
                b1043 := true;
                b1045 := true;
                b1047 := true;
                b1049 := true;
                b1051 := true;
                b1053 := true;
                b1055 := true;
                b1057 := true;
                b1059 := true;
                b1061 := true;
                null;
                null;
                -- got x0@225 in r999
                -- got x1@226 in r1001
                -- got x2@227 in r1003
                -- got x3@228 in r1005
                -- got w1'@223 in r988
                -- got w2'@224 in r990
                -- got x6@22B in r1011
                -- got x7@22C in r1013
                -- got x8@22D in r1015
                -- got x9@22E in r1017
                -- got xa@22F in r1019
                -- got xb@22G in r1021
                -- got xc@22H in r1023
                -- got xd@22I in r1025
                -- got xe@22J in r1027
                -- got xf@22K in r1029
                r1064 := (r999 & r1001 & r1003 & r1005 & r988 & r990 & r1011 & r1013 & r1015 & r1017 & r1019 & r1021 & r1023 & r1025 & r1027 & r1029);
                r986 := r1064;
                -- end case
                statevar1 := r986;
                r1086 := "1";
                r1089 := "0000000000000000000000000000000000000000000000000000000000000000";
                r1088 := (r1086 & r1089);
                output_tmp := r1088;
                control := STATE1094;
                goto_L7852 := true;
              end if;
              goto_L7852 := goto_L7852;
            end if;
            goto_L7852 := goto_L7852;
            if (NOT goto_L7852) then
              null; -- label L842
              r841 := statevar1;
              null;
              null;
              -- got w1@219 in r831
              -- got w2@21A in r833
              -- got hw@21B in r841
              r844 := (r831 & r833 & r841);
              -- final pat
              r852 := r844(0 to 31);
              r854 := r844(32 to 63);
              r856 := r844(64 to 575);
              b858 := true;
              b860 := true;
              -- final pat
              r863 := r856(0 to 31);
              r865 := r856(32 to 63);
              r867 := r856(64 to 95);
              r869 := r856(96 to 127);
              r871 := r856(128 to 159);
              r873 := r856(160 to 191);
              r875 := r856(192 to 223);
              r877 := r856(224 to 255);
              r879 := r856(256 to 287);
              r881 := r856(288 to 319);
              r883 := r856(320 to 351);
              r885 := r856(352 to 383);
              r887 := r856(384 to 415);
              r889 := r856(416 to 447);
              r891 := r856(448 to 479);
              r893 := r856(480 to 511);
              b895 := true;
              b897 := true;
              b899 := true;
              b901 := true;
              b903 := true;
              b905 := true;
              b907 := true;
              b909 := true;
              b911 := true;
              b913 := true;
              b915 := true;
              b917 := true;
              b919 := true;
              b921 := true;
              b923 := true;
              b925 := true;
              null;
              null;
              -- got x0@21E in r863
              -- got x1@21F in r865
              -- got w1'@21C in r852
              -- got w2'@21D in r854
              -- got x4@21I in r871
              -- got x5@21J in r873
              -- got x6@21K in r875
              -- got x7@21L in r877
              -- got x8@21M in r879
              -- got x9@21N in r881
              -- got xa@21O in r883
              -- got xb@21P in r885
              -- got xc@21Q in r887
              -- got xd@21R in r889
              -- got xe@21S in r891
              -- got xf@21T in r893
              r928 := (r863 & r865 & r852 & r854 & r871 & r873 & r875 & r877 & r879 & r881 & r883 & r885 & r887 & r889 & r891 & r893);
              r850 := r928;
              -- end case
              statevar1 := r850;
              r950 := "1";
              r953 := "0000000000000000000000000000000000000000000000000000000000000000";
              r952 := (r950 & r953);
              output_tmp := r952;
              control := STATE958;
              goto_L7852 := true;
            end if;
            goto_L7852 := goto_L7852;
          end if;
          goto_L7852 := goto_L7852;
          if (NOT goto_L7852) then
            null; -- label L706
            r705 := statevar1;
            null;
            null;
            -- got w1@20I in r695
            -- got w2@20J in r697
            -- got hw@20K in r705
            r708 := (r695 & r697 & r705);
            -- final pat
            r716 := r708(0 to 31);
            r718 := r708(32 to 63);
            r720 := r708(64 to 575);
            b722 := true;
            b724 := true;
            -- final pat
            r727 := r720(0 to 31);
            r729 := r720(32 to 63);
            r731 := r720(64 to 95);
            r733 := r720(96 to 127);
            r735 := r720(128 to 159);
            r737 := r720(160 to 191);
            r739 := r720(192 to 223);
            r741 := r720(224 to 255);
            r743 := r720(256 to 287);
            r745 := r720(288 to 319);
            r747 := r720(320 to 351);
            r749 := r720(352 to 383);
            r751 := r720(384 to 415);
            r753 := r720(416 to 447);
            r755 := r720(448 to 479);
            r757 := r720(480 to 511);
            b759 := true;
            b761 := true;
            b763 := true;
            b765 := true;
            b767 := true;
            b769 := true;
            b771 := true;
            b773 := true;
            b775 := true;
            b777 := true;
            b779 := true;
            b781 := true;
            b783 := true;
            b785 := true;
            b787 := true;
            b789 := true;
            null;
            null;
            -- got w1'@20L in r716
            -- got w2'@20M in r718
            -- got x2@20P in r731
            -- got x3@20Q in r733
            -- got x4@20R in r735
            -- got x5@20S in r737
            -- got x6@20T in r739
            -- got x7@20U in r741
            -- got x8@20V in r743
            -- got x9@210 in r745
            -- got xa@211 in r747
            -- got xb@212 in r749
            -- got xc@213 in r751
            -- got xd@214 in r753
            -- got xe@215 in r755
            -- got xf@216 in r757
            r792 := (r716 & r718 & r731 & r733 & r735 & r737 & r739 & r741 & r743 & r745 & r747 & r749 & r751 & r753 & r755 & r757);
            r714 := r792;
            -- end case
            statevar1 := r714;
            r814 := "1";
            r817 := "0000000000000000000000000000000000000000000000000000000000000000";
            r816 := (r814 & r817);
            output_tmp := r816;
            control := STATE822;
            goto_L7852 := true;
          end if;
          goto_L7852 := goto_L7852;
        end if;
        goto_L7852 := goto_L7852;
        if (NOT goto_L7852) then
          null; -- label L567
          r566 := rewire_MaininitialSHA256State_28;
          statevar2 := r566;
          r569 := statevar1;
          null;
          null;
          -- got w1@1VQ in r18
          -- got w2@1VR in r20
          -- got hw@1VT in r569
          r572 := (r18 & r20 & r569);
          -- final pat
          r580 := r572(0 to 31);
          r582 := r572(32 to 63);
          r584 := r572(64 to 575);
          b586 := true;
          b588 := true;
          -- final pat
          r591 := r584(0 to 31);
          r593 := r584(32 to 63);
          r595 := r584(64 to 95);
          r597 := r584(96 to 127);
          r599 := r584(128 to 159);
          r601 := r584(160 to 191);
          r603 := r584(192 to 223);
          r605 := r584(224 to 255);
          r607 := r584(256 to 287);
          r609 := r584(288 to 319);
          r611 := r584(320 to 351);
          r613 := r584(352 to 383);
          r615 := r584(384 to 415);
          r617 := r584(416 to 447);
          r619 := r584(448 to 479);
          r621 := r584(480 to 511);
          b623 := true;
          b625 := true;
          b627 := true;
          b629 := true;
          b631 := true;
          b633 := true;
          b635 := true;
          b637 := true;
          b639 := true;
          b641 := true;
          b643 := true;
          b645 := true;
          b647 := true;
          b649 := true;
          b651 := true;
          b653 := true;
          null;
          null;
          -- got w1'@1VU in r580
          -- got w2'@1VV in r582
          -- got x2@202 in r595
          -- got x3@203 in r597
          -- got x4@204 in r599
          -- got x5@205 in r601
          -- got x6@206 in r603
          -- got x7@207 in r605
          -- got x8@208 in r607
          -- got x9@209 in r609
          -- got xa@20A in r611
          -- got xb@20B in r613
          -- got xc@20C in r615
          -- got xd@20D in r617
          -- got xe@20E in r619
          -- got xf@20F in r621
          r656 := (r580 & r582 & r595 & r597 & r599 & r601 & r603 & r605 & r607 & r609 & r611 & r613 & r615 & r617 & r619 & r621);
          r578 := r656;
          -- end case
          statevar1 := r578;
          r678 := "1";
          r681 := "0000000000000000000000000000000000000000000000000000000000000000";
          r680 := (r678 & r681);
          output_tmp := r680;
          control := STATE686;
          goto_L7852 := true;
        end if;
        goto_L7852 := goto_L7852;
      end if;
      goto_L7852 := goto_L7852;
    end if;
    goto_L7852 := goto_L7852;
    if (NOT goto_L7852) then
      null; -- label L0
      -- START
      -- Maindevsha256' in
      r3 := "1";
      r6 := "0000000000000000000000000000000000000000000000000000000000000000";
      r5 := (r3 & r6);
      output_tmp := r5;
      control := STATE11;
      goto_L7852 := true;
    end if;
    goto_L7852 := goto_L7852;
    null; -- label L7852
    -- EXIT
    -- Write back reg temps.
    control_flop_next <= control;
    goto_L7851_flop_next <= goto_L7851;
    goto_L7844_flop_next <= goto_L7844;
    goto_L7806_flop_next <= goto_L7806;
    goto_L7767_flop_next <= goto_L7767;
    goto_L7728_flop_next <= goto_L7728;
    goto_L7570_flop_next <= goto_L7570;
    goto_L7690_flop_next <= goto_L7690;
    goto_L7575_flop_next <= goto_L7575;
    goto_L1784_flop_next <= goto_L1784;
    goto_L1785_flop_next <= goto_L1785;
    goto_L1638_flop_next <= goto_L1638;
    goto_L1502_flop_next <= goto_L1502;
    goto_L1366_flop_next <= goto_L1366;
    goto_L1230_flop_next <= goto_L1230;
    goto_L1094_flop_next <= goto_L1094;
    goto_L958_flop_next <= goto_L958;
    goto_L822_flop_next <= goto_L822;
    goto_L686_flop_next <= goto_L686;
    goto_L11_flop_next <= goto_L11;
    goto_L13_flop_next <= goto_L13;
    goto_L690_flop_next <= goto_L690;
    goto_L826_flop_next <= goto_L826;
    goto_L962_flop_next <= goto_L962;
    goto_L1098_flop_next <= goto_L1098;
    goto_L1234_flop_next <= goto_L1234;
    goto_L1370_flop_next <= goto_L1370;
    goto_L1506_flop_next <= goto_L1506;
    goto_L1642_flop_next <= goto_L1642;
    goto_L7693_flop_next <= goto_L7693;
    goto_L7732_flop_next <= goto_L7732;
    goto_L7771_flop_next <= goto_L7771;
    goto_L7810_flop_next <= goto_L7810;
    goto_L7777_flop_next <= goto_L7777;
    goto_L7738_flop_next <= goto_L7738;
    goto_L7699_flop_next <= goto_L7699;
    goto_L1658_flop_next <= goto_L1658;
    goto_L1522_flop_next <= goto_L1522;
    goto_L1386_flop_next <= goto_L1386;
    goto_L1250_flop_next <= goto_L1250;
    goto_L1114_flop_next <= goto_L1114;
    goto_L978_flop_next <= goto_L978;
    goto_L842_flop_next <= goto_L842;
    goto_L706_flop_next <= goto_L706;
    goto_L567_flop_next <= goto_L567;
    goto_L0_flop_next <= goto_L0;
    goto_L7852_flop_next <= goto_L7852;
    r7843_flop_next <= r7843;
    r7840_flop_next <= r7840;
    r7817_flop_next <= r7817;
    r7814_flop_next <= r7814;
    r7805_flop_next <= r7805;
    r7802_flop_next <= r7802;
    r7779_flop_next <= r7779;
    r7776_flop_next <= r7776;
    b7774_flop_next <= b7774;
    r7766_flop_next <= r7766;
    r7763_flop_next <= r7763;
    r7740_flop_next <= r7740;
    r7737_flop_next <= r7737;
    b7735_flop_next <= b7735;
    r7727_flop_next <= r7727;
    r7724_flop_next <= r7724;
    r7701_flop_next <= r7701;
    r7698_flop_next <= r7698;
    b7696_flop_next <= b7696;
    r7679_flop_next <= r7679;
    r7675_flop_next <= r7675;
    r7671_flop_next <= r7671;
    r7667_flop_next <= r7667;
    r7663_flop_next <= r7663;
    r7659_flop_next <= r7659;
    r7655_flop_next <= r7655;
    r7651_flop_next <= r7651;
    r7647_flop_next <= r7647;
    b7644_flop_next <= b7644;
    b7642_flop_next <= b7642;
    b7640_flop_next <= b7640;
    b7638_flop_next <= b7638;
    b7636_flop_next <= b7636;
    b7634_flop_next <= b7634;
    b7632_flop_next <= b7632;
    b7630_flop_next <= b7630;
    r7628_flop_next <= r7628;
    r7626_flop_next <= r7626;
    r7624_flop_next <= r7624;
    r7622_flop_next <= r7622;
    r7620_flop_next <= r7620;
    r7618_flop_next <= r7618;
    r7616_flop_next <= r7616;
    r7614_flop_next <= r7614;
    r7610_flop_next <= r7610;
    b7608_flop_next <= b7608;
    b7606_flop_next <= b7606;
    b7604_flop_next <= b7604;
    b7602_flop_next <= b7602;
    b7600_flop_next <= b7600;
    b7598_flop_next <= b7598;
    b7596_flop_next <= b7596;
    b7594_flop_next <= b7594;
    r7592_flop_next <= r7592;
    r7590_flop_next <= r7590;
    r7588_flop_next <= r7588;
    r7586_flop_next <= r7586;
    r7584_flop_next <= r7584;
    r7582_flop_next <= r7582;
    r7580_flop_next <= r7580;
    r7578_flop_next <= r7578;
    r7574_flop_next <= r7574;
    b7572_flop_next <= b7572;
    r7569_flop_next <= r7569;
    r7565_flop_next <= r7565;
    r7564_flop_next <= r7564;
    r7562_flop_next <= r7562;
    r7558_flop_next <= r7558;
    r7300_flop_next <= r7300;
    r7296_flop_next <= r7296;
    r7292_flop_next <= r7292;
    r2874_flop_next <= r2874;
    r2376_flop_next <= r2376;
    r2375_flop_next <= r2375;
    r2374_flop_next <= r2374;
    r2371_flop_next <= r2371;
    r2365_flop_next <= r2365;
    r1862_flop_next <= r1862;
    b1859_flop_next <= b1859;
    b1857_flop_next <= b1857;
    b1855_flop_next <= b1855;
    b1853_flop_next <= b1853;
    b1851_flop_next <= b1851;
    b1849_flop_next <= b1849;
    b1847_flop_next <= b1847;
    b1845_flop_next <= b1845;
    b1843_flop_next <= b1843;
    b1841_flop_next <= b1841;
    b1839_flop_next <= b1839;
    b1837_flop_next <= b1837;
    b1835_flop_next <= b1835;
    b1833_flop_next <= b1833;
    b1831_flop_next <= b1831;
    b1829_flop_next <= b1829;
    r1827_flop_next <= r1827;
    r1825_flop_next <= r1825;
    r1823_flop_next <= r1823;
    r1821_flop_next <= r1821;
    r1819_flop_next <= r1819;
    r1817_flop_next <= r1817;
    r1815_flop_next <= r1815;
    r1813_flop_next <= r1813;
    r1811_flop_next <= r1811;
    r1809_flop_next <= r1809;
    r1807_flop_next <= r1807;
    r1805_flop_next <= r1805;
    r1803_flop_next <= r1803;
    r1801_flop_next <= r1801;
    r1799_flop_next <= r1799;
    r1797_flop_next <= r1797;
    r1795_flop_next <= r1795;
    r1792_flop_next <= r1792;
    r1790_flop_next <= r1790;
    r1787_flop_next <= r1787;
    r1783_flop_next <= r1783;
    r1779_flop_next <= r1779;
    r1778_flop_next <= r1778;
    r1776_flop_next <= r1776;
    r1754_flop_next <= r1754;
    b1751_flop_next <= b1751;
    b1749_flop_next <= b1749;
    b1747_flop_next <= b1747;
    b1745_flop_next <= b1745;
    b1743_flop_next <= b1743;
    b1741_flop_next <= b1741;
    b1739_flop_next <= b1739;
    b1737_flop_next <= b1737;
    b1735_flop_next <= b1735;
    b1733_flop_next <= b1733;
    b1731_flop_next <= b1731;
    b1729_flop_next <= b1729;
    b1727_flop_next <= b1727;
    b1725_flop_next <= b1725;
    b1723_flop_next <= b1723;
    b1721_flop_next <= b1721;
    r1719_flop_next <= r1719;
    r1717_flop_next <= r1717;
    r1715_flop_next <= r1715;
    r1713_flop_next <= r1713;
    r1711_flop_next <= r1711;
    r1709_flop_next <= r1709;
    r1707_flop_next <= r1707;
    r1705_flop_next <= r1705;
    r1703_flop_next <= r1703;
    r1701_flop_next <= r1701;
    r1699_flop_next <= r1699;
    r1697_flop_next <= r1697;
    r1695_flop_next <= r1695;
    r1693_flop_next <= r1693;
    r1691_flop_next <= r1691;
    r1689_flop_next <= r1689;
    b1686_flop_next <= b1686;
    b1684_flop_next <= b1684;
    r1682_flop_next <= r1682;
    r1680_flop_next <= r1680;
    r1678_flop_next <= r1678;
    r1676_flop_next <= r1676;
    r1670_flop_next <= r1670;
    r1667_flop_next <= r1667;
    r1663_flop_next <= r1663;
    r1659_flop_next <= r1659;
    r1657_flop_next <= r1657;
    b1655_flop_next <= b1655;
    b1653_flop_next <= b1653;
    b1651_flop_next <= b1651;
    r1649_flop_next <= r1649;
    r1647_flop_next <= r1647;
    b1645_flop_next <= b1645;
    r1637_flop_next <= r1637;
    r1633_flop_next <= r1633;
    r1632_flop_next <= r1632;
    r1630_flop_next <= r1630;
    r1608_flop_next <= r1608;
    b1605_flop_next <= b1605;
    b1603_flop_next <= b1603;
    b1601_flop_next <= b1601;
    b1599_flop_next <= b1599;
    b1597_flop_next <= b1597;
    b1595_flop_next <= b1595;
    b1593_flop_next <= b1593;
    b1591_flop_next <= b1591;
    b1589_flop_next <= b1589;
    b1587_flop_next <= b1587;
    b1585_flop_next <= b1585;
    b1583_flop_next <= b1583;
    b1581_flop_next <= b1581;
    b1579_flop_next <= b1579;
    b1577_flop_next <= b1577;
    b1575_flop_next <= b1575;
    r1573_flop_next <= r1573;
    r1571_flop_next <= r1571;
    r1569_flop_next <= r1569;
    r1567_flop_next <= r1567;
    r1565_flop_next <= r1565;
    r1563_flop_next <= r1563;
    r1561_flop_next <= r1561;
    r1559_flop_next <= r1559;
    r1557_flop_next <= r1557;
    r1555_flop_next <= r1555;
    r1553_flop_next <= r1553;
    r1551_flop_next <= r1551;
    r1549_flop_next <= r1549;
    r1547_flop_next <= r1547;
    r1545_flop_next <= r1545;
    r1543_flop_next <= r1543;
    b1540_flop_next <= b1540;
    b1538_flop_next <= b1538;
    r1536_flop_next <= r1536;
    r1534_flop_next <= r1534;
    r1532_flop_next <= r1532;
    r1530_flop_next <= r1530;
    r1524_flop_next <= r1524;
    r1521_flop_next <= r1521;
    b1519_flop_next <= b1519;
    b1517_flop_next <= b1517;
    b1515_flop_next <= b1515;
    r1513_flop_next <= r1513;
    r1511_flop_next <= r1511;
    b1509_flop_next <= b1509;
    r1501_flop_next <= r1501;
    r1497_flop_next <= r1497;
    r1496_flop_next <= r1496;
    r1494_flop_next <= r1494;
    r1472_flop_next <= r1472;
    b1469_flop_next <= b1469;
    b1467_flop_next <= b1467;
    b1465_flop_next <= b1465;
    b1463_flop_next <= b1463;
    b1461_flop_next <= b1461;
    b1459_flop_next <= b1459;
    b1457_flop_next <= b1457;
    b1455_flop_next <= b1455;
    b1453_flop_next <= b1453;
    b1451_flop_next <= b1451;
    b1449_flop_next <= b1449;
    b1447_flop_next <= b1447;
    b1445_flop_next <= b1445;
    b1443_flop_next <= b1443;
    b1441_flop_next <= b1441;
    b1439_flop_next <= b1439;
    r1437_flop_next <= r1437;
    r1435_flop_next <= r1435;
    r1433_flop_next <= r1433;
    r1431_flop_next <= r1431;
    r1429_flop_next <= r1429;
    r1427_flop_next <= r1427;
    r1425_flop_next <= r1425;
    r1423_flop_next <= r1423;
    r1421_flop_next <= r1421;
    r1419_flop_next <= r1419;
    r1417_flop_next <= r1417;
    r1415_flop_next <= r1415;
    r1413_flop_next <= r1413;
    r1411_flop_next <= r1411;
    r1409_flop_next <= r1409;
    r1407_flop_next <= r1407;
    b1404_flop_next <= b1404;
    b1402_flop_next <= b1402;
    r1400_flop_next <= r1400;
    r1398_flop_next <= r1398;
    r1396_flop_next <= r1396;
    r1394_flop_next <= r1394;
    r1388_flop_next <= r1388;
    r1385_flop_next <= r1385;
    b1383_flop_next <= b1383;
    b1381_flop_next <= b1381;
    b1379_flop_next <= b1379;
    r1377_flop_next <= r1377;
    r1375_flop_next <= r1375;
    b1373_flop_next <= b1373;
    r1365_flop_next <= r1365;
    r1361_flop_next <= r1361;
    r1360_flop_next <= r1360;
    r1358_flop_next <= r1358;
    r1336_flop_next <= r1336;
    b1333_flop_next <= b1333;
    b1331_flop_next <= b1331;
    b1329_flop_next <= b1329;
    b1327_flop_next <= b1327;
    b1325_flop_next <= b1325;
    b1323_flop_next <= b1323;
    b1321_flop_next <= b1321;
    b1319_flop_next <= b1319;
    b1317_flop_next <= b1317;
    b1315_flop_next <= b1315;
    b1313_flop_next <= b1313;
    b1311_flop_next <= b1311;
    b1309_flop_next <= b1309;
    b1307_flop_next <= b1307;
    b1305_flop_next <= b1305;
    b1303_flop_next <= b1303;
    r1301_flop_next <= r1301;
    r1299_flop_next <= r1299;
    r1297_flop_next <= r1297;
    r1295_flop_next <= r1295;
    r1293_flop_next <= r1293;
    r1291_flop_next <= r1291;
    r1289_flop_next <= r1289;
    r1287_flop_next <= r1287;
    r1285_flop_next <= r1285;
    r1283_flop_next <= r1283;
    r1281_flop_next <= r1281;
    r1279_flop_next <= r1279;
    r1277_flop_next <= r1277;
    r1275_flop_next <= r1275;
    r1273_flop_next <= r1273;
    r1271_flop_next <= r1271;
    b1268_flop_next <= b1268;
    b1266_flop_next <= b1266;
    r1264_flop_next <= r1264;
    r1262_flop_next <= r1262;
    r1260_flop_next <= r1260;
    r1258_flop_next <= r1258;
    r1252_flop_next <= r1252;
    r1249_flop_next <= r1249;
    b1247_flop_next <= b1247;
    b1245_flop_next <= b1245;
    b1243_flop_next <= b1243;
    r1241_flop_next <= r1241;
    r1239_flop_next <= r1239;
    b1237_flop_next <= b1237;
    r1229_flop_next <= r1229;
    r1225_flop_next <= r1225;
    r1224_flop_next <= r1224;
    r1222_flop_next <= r1222;
    r1200_flop_next <= r1200;
    b1197_flop_next <= b1197;
    b1195_flop_next <= b1195;
    b1193_flop_next <= b1193;
    b1191_flop_next <= b1191;
    b1189_flop_next <= b1189;
    b1187_flop_next <= b1187;
    b1185_flop_next <= b1185;
    b1183_flop_next <= b1183;
    b1181_flop_next <= b1181;
    b1179_flop_next <= b1179;
    b1177_flop_next <= b1177;
    b1175_flop_next <= b1175;
    b1173_flop_next <= b1173;
    b1171_flop_next <= b1171;
    b1169_flop_next <= b1169;
    b1167_flop_next <= b1167;
    r1165_flop_next <= r1165;
    r1163_flop_next <= r1163;
    r1161_flop_next <= r1161;
    r1159_flop_next <= r1159;
    r1157_flop_next <= r1157;
    r1155_flop_next <= r1155;
    r1153_flop_next <= r1153;
    r1151_flop_next <= r1151;
    r1149_flop_next <= r1149;
    r1147_flop_next <= r1147;
    r1145_flop_next <= r1145;
    r1143_flop_next <= r1143;
    r1141_flop_next <= r1141;
    r1139_flop_next <= r1139;
    r1137_flop_next <= r1137;
    r1135_flop_next <= r1135;
    b1132_flop_next <= b1132;
    b1130_flop_next <= b1130;
    r1128_flop_next <= r1128;
    r1126_flop_next <= r1126;
    r1124_flop_next <= r1124;
    r1122_flop_next <= r1122;
    r1116_flop_next <= r1116;
    r1113_flop_next <= r1113;
    b1111_flop_next <= b1111;
    b1109_flop_next <= b1109;
    b1107_flop_next <= b1107;
    r1105_flop_next <= r1105;
    r1103_flop_next <= r1103;
    b1101_flop_next <= b1101;
    r1093_flop_next <= r1093;
    r1089_flop_next <= r1089;
    r1088_flop_next <= r1088;
    r1086_flop_next <= r1086;
    r1064_flop_next <= r1064;
    b1061_flop_next <= b1061;
    b1059_flop_next <= b1059;
    b1057_flop_next <= b1057;
    b1055_flop_next <= b1055;
    b1053_flop_next <= b1053;
    b1051_flop_next <= b1051;
    b1049_flop_next <= b1049;
    b1047_flop_next <= b1047;
    b1045_flop_next <= b1045;
    b1043_flop_next <= b1043;
    b1041_flop_next <= b1041;
    b1039_flop_next <= b1039;
    b1037_flop_next <= b1037;
    b1035_flop_next <= b1035;
    b1033_flop_next <= b1033;
    b1031_flop_next <= b1031;
    r1029_flop_next <= r1029;
    r1027_flop_next <= r1027;
    r1025_flop_next <= r1025;
    r1023_flop_next <= r1023;
    r1021_flop_next <= r1021;
    r1019_flop_next <= r1019;
    r1017_flop_next <= r1017;
    r1015_flop_next <= r1015;
    r1013_flop_next <= r1013;
    r1011_flop_next <= r1011;
    r1009_flop_next <= r1009;
    r1007_flop_next <= r1007;
    r1005_flop_next <= r1005;
    r1003_flop_next <= r1003;
    r1001_flop_next <= r1001;
    r999_flop_next <= r999;
    b996_flop_next <= b996;
    b994_flop_next <= b994;
    r992_flop_next <= r992;
    r990_flop_next <= r990;
    r988_flop_next <= r988;
    r986_flop_next <= r986;
    r980_flop_next <= r980;
    r977_flop_next <= r977;
    b975_flop_next <= b975;
    b973_flop_next <= b973;
    b971_flop_next <= b971;
    r969_flop_next <= r969;
    r967_flop_next <= r967;
    b965_flop_next <= b965;
    r957_flop_next <= r957;
    r953_flop_next <= r953;
    r952_flop_next <= r952;
    r950_flop_next <= r950;
    r928_flop_next <= r928;
    b925_flop_next <= b925;
    b923_flop_next <= b923;
    b921_flop_next <= b921;
    b919_flop_next <= b919;
    b917_flop_next <= b917;
    b915_flop_next <= b915;
    b913_flop_next <= b913;
    b911_flop_next <= b911;
    b909_flop_next <= b909;
    b907_flop_next <= b907;
    b905_flop_next <= b905;
    b903_flop_next <= b903;
    b901_flop_next <= b901;
    b899_flop_next <= b899;
    b897_flop_next <= b897;
    b895_flop_next <= b895;
    r893_flop_next <= r893;
    r891_flop_next <= r891;
    r889_flop_next <= r889;
    r887_flop_next <= r887;
    r885_flop_next <= r885;
    r883_flop_next <= r883;
    r881_flop_next <= r881;
    r879_flop_next <= r879;
    r877_flop_next <= r877;
    r875_flop_next <= r875;
    r873_flop_next <= r873;
    r871_flop_next <= r871;
    r869_flop_next <= r869;
    r867_flop_next <= r867;
    r865_flop_next <= r865;
    r863_flop_next <= r863;
    b860_flop_next <= b860;
    b858_flop_next <= b858;
    r856_flop_next <= r856;
    r854_flop_next <= r854;
    r852_flop_next <= r852;
    r850_flop_next <= r850;
    r844_flop_next <= r844;
    r841_flop_next <= r841;
    b839_flop_next <= b839;
    b837_flop_next <= b837;
    b835_flop_next <= b835;
    r833_flop_next <= r833;
    r831_flop_next <= r831;
    b829_flop_next <= b829;
    r821_flop_next <= r821;
    r817_flop_next <= r817;
    r816_flop_next <= r816;
    r814_flop_next <= r814;
    r792_flop_next <= r792;
    b789_flop_next <= b789;
    b787_flop_next <= b787;
    b785_flop_next <= b785;
    b783_flop_next <= b783;
    b781_flop_next <= b781;
    b779_flop_next <= b779;
    b777_flop_next <= b777;
    b775_flop_next <= b775;
    b773_flop_next <= b773;
    b771_flop_next <= b771;
    b769_flop_next <= b769;
    b767_flop_next <= b767;
    b765_flop_next <= b765;
    b763_flop_next <= b763;
    b761_flop_next <= b761;
    b759_flop_next <= b759;
    r757_flop_next <= r757;
    r755_flop_next <= r755;
    r753_flop_next <= r753;
    r751_flop_next <= r751;
    r749_flop_next <= r749;
    r747_flop_next <= r747;
    r745_flop_next <= r745;
    r743_flop_next <= r743;
    r741_flop_next <= r741;
    r739_flop_next <= r739;
    r737_flop_next <= r737;
    r735_flop_next <= r735;
    r733_flop_next <= r733;
    r731_flop_next <= r731;
    r729_flop_next <= r729;
    r727_flop_next <= r727;
    b724_flop_next <= b724;
    b722_flop_next <= b722;
    r720_flop_next <= r720;
    r718_flop_next <= r718;
    r716_flop_next <= r716;
    r714_flop_next <= r714;
    r708_flop_next <= r708;
    r705_flop_next <= r705;
    b703_flop_next <= b703;
    b701_flop_next <= b701;
    b699_flop_next <= b699;
    r697_flop_next <= r697;
    r695_flop_next <= r695;
    b693_flop_next <= b693;
    r685_flop_next <= r685;
    r681_flop_next <= r681;
    r680_flop_next <= r680;
    r678_flop_next <= r678;
    r656_flop_next <= r656;
    b653_flop_next <= b653;
    b651_flop_next <= b651;
    b649_flop_next <= b649;
    b647_flop_next <= b647;
    b645_flop_next <= b645;
    b643_flop_next <= b643;
    b641_flop_next <= b641;
    b639_flop_next <= b639;
    b637_flop_next <= b637;
    b635_flop_next <= b635;
    b633_flop_next <= b633;
    b631_flop_next <= b631;
    b629_flop_next <= b629;
    b627_flop_next <= b627;
    b625_flop_next <= b625;
    b623_flop_next <= b623;
    r621_flop_next <= r621;
    r619_flop_next <= r619;
    r617_flop_next <= r617;
    r615_flop_next <= r615;
    r613_flop_next <= r613;
    r611_flop_next <= r611;
    r609_flop_next <= r609;
    r607_flop_next <= r607;
    r605_flop_next <= r605;
    r603_flop_next <= r603;
    r601_flop_next <= r601;
    r599_flop_next <= r599;
    r597_flop_next <= r597;
    r595_flop_next <= r595;
    r593_flop_next <= r593;
    r591_flop_next <= r591;
    b588_flop_next <= b588;
    b586_flop_next <= b586;
    r584_flop_next <= r584;
    r582_flop_next <= r582;
    r580_flop_next <= r580;
    r578_flop_next <= r578;
    r572_flop_next <= r572;
    r569_flop_next <= r569;
    r566_flop_next <= r566;
    b26_flop_next <= b26;
    b24_flop_next <= b24;
    b22_flop_next <= b22;
    r20_flop_next <= r20;
    r18_flop_next <= r18;
    b16_flop_next <= b16;
    r12_flop_next <= r12;
    r10_flop_next <= r10;
    r6_flop_next <= r6;
    r5_flop_next <= r5;
    r3_flop_next <= r3;
    statevar0_flop_next <= statevar0;
    statevar1_flop_next <= statevar1;
    statevar2_flop_next <= statevar2;
    statevar3_flop_next <= statevar3;
    -- Update output line.
    output <= output_tmp;
  end process;

  -- Flip flop update process.
  process (clk,input,goto_L7851_flop_next,goto_L7844_flop_next,goto_L7806_flop_next,goto_L7767_flop_next,goto_L7728_flop_next,goto_L7570_flop_next,goto_L7690_flop_next,goto_L7575_flop_next,goto_L1784_flop_next,goto_L1785_flop_next,goto_L1638_flop_next,goto_L1502_flop_next,goto_L1366_flop_next,goto_L1230_flop_next,goto_L1094_flop_next,goto_L958_flop_next,goto_L822_flop_next,goto_L686_flop_next,goto_L11_flop_next,goto_L13_flop_next,goto_L690_flop_next,goto_L826_flop_next,goto_L962_flop_next,goto_L1098_flop_next,goto_L1234_flop_next,goto_L1370_flop_next,goto_L1506_flop_next,goto_L1642_flop_next,goto_L7693_flop_next,goto_L7732_flop_next,goto_L7771_flop_next,goto_L7810_flop_next,goto_L7777_flop_next,goto_L7738_flop_next,goto_L7699_flop_next,goto_L1658_flop_next,goto_L1522_flop_next,goto_L1386_flop_next,goto_L1250_flop_next,goto_L1114_flop_next,goto_L978_flop_next,goto_L842_flop_next,goto_L706_flop_next,goto_L567_flop_next,goto_L0_flop_next,goto_L7852_flop_next,r7843_flop_next,r7840_flop_next,r7817_flop_next,r7814_flop_next,r7805_flop_next,r7802_flop_next,r7779_flop_next,r7776_flop_next,b7774_flop_next,r7766_flop_next,r7763_flop_next,r7740_flop_next,r7737_flop_next,b7735_flop_next,r7727_flop_next,r7724_flop_next,r7701_flop_next,r7698_flop_next,b7696_flop_next,r7679_flop_next,r7675_flop_next,r7671_flop_next,r7667_flop_next,r7663_flop_next,r7659_flop_next,r7655_flop_next,r7651_flop_next,r7647_flop_next,b7644_flop_next,b7642_flop_next,b7640_flop_next,b7638_flop_next,b7636_flop_next,b7634_flop_next,b7632_flop_next,b7630_flop_next,r7628_flop_next,r7626_flop_next,r7624_flop_next,r7622_flop_next,r7620_flop_next,r7618_flop_next,r7616_flop_next,r7614_flop_next,r7610_flop_next,b7608_flop_next,b7606_flop_next,b7604_flop_next,b7602_flop_next,b7600_flop_next,b7598_flop_next,b7596_flop_next,b7594_flop_next,r7592_flop_next,r7590_flop_next,r7588_flop_next,r7586_flop_next,r7584_flop_next,r7582_flop_next,r7580_flop_next,r7578_flop_next,r7574_flop_next,b7572_flop_next,r7569_flop_next,r7565_flop_next,r7564_flop_next,r7562_flop_next,r7558_flop_next,r7300_flop_next,r7296_flop_next,r7292_flop_next,r2874_flop_next,r2376_flop_next,r2375_flop_next,r2374_flop_next,r2371_flop_next,r2365_flop_next,r1862_flop_next,b1859_flop_next,b1857_flop_next,b1855_flop_next,b1853_flop_next,b1851_flop_next,b1849_flop_next,b1847_flop_next,b1845_flop_next,b1843_flop_next,b1841_flop_next,b1839_flop_next,b1837_flop_next,b1835_flop_next,b1833_flop_next,b1831_flop_next,b1829_flop_next,r1827_flop_next,r1825_flop_next,r1823_flop_next,r1821_flop_next,r1819_flop_next,r1817_flop_next,r1815_flop_next,r1813_flop_next,r1811_flop_next,r1809_flop_next,r1807_flop_next,r1805_flop_next,r1803_flop_next,r1801_flop_next,r1799_flop_next,r1797_flop_next,r1795_flop_next,r1792_flop_next,r1790_flop_next,r1787_flop_next,r1783_flop_next,r1779_flop_next,r1778_flop_next,r1776_flop_next,r1754_flop_next,b1751_flop_next,b1749_flop_next,b1747_flop_next,b1745_flop_next,b1743_flop_next,b1741_flop_next,b1739_flop_next,b1737_flop_next,b1735_flop_next,b1733_flop_next,b1731_flop_next,b1729_flop_next,b1727_flop_next,b1725_flop_next,b1723_flop_next,b1721_flop_next,r1719_flop_next,r1717_flop_next,r1715_flop_next,r1713_flop_next,r1711_flop_next,r1709_flop_next,r1707_flop_next,r1705_flop_next,r1703_flop_next,r1701_flop_next,r1699_flop_next,r1697_flop_next,r1695_flop_next,r1693_flop_next,r1691_flop_next,r1689_flop_next,b1686_flop_next,b1684_flop_next,r1682_flop_next,r1680_flop_next,r1678_flop_next,r1676_flop_next,r1670_flop_next,r1667_flop_next,r1663_flop_next,r1659_flop_next,r1657_flop_next,b1655_flop_next,b1653_flop_next,b1651_flop_next,r1649_flop_next,r1647_flop_next,b1645_flop_next,r1637_flop_next,r1633_flop_next,r1632_flop_next,r1630_flop_next,r1608_flop_next,b1605_flop_next,b1603_flop_next,b1601_flop_next,b1599_flop_next,b1597_flop_next,b1595_flop_next,b1593_flop_next,b1591_flop_next,b1589_flop_next,b1587_flop_next,b1585_flop_next,b1583_flop_next,b1581_flop_next,b1579_flop_next,b1577_flop_next,b1575_flop_next,r1573_flop_next,r1571_flop_next,r1569_flop_next,r1567_flop_next,r1565_flop_next,r1563_flop_next,r1561_flop_next,r1559_flop_next,r1557_flop_next,r1555_flop_next,r1553_flop_next,r1551_flop_next,r1549_flop_next,r1547_flop_next,r1545_flop_next,r1543_flop_next,b1540_flop_next,b1538_flop_next,r1536_flop_next,r1534_flop_next,r1532_flop_next,r1530_flop_next,r1524_flop_next,r1521_flop_next,b1519_flop_next,b1517_flop_next,b1515_flop_next,r1513_flop_next,r1511_flop_next,b1509_flop_next,r1501_flop_next,r1497_flop_next,r1496_flop_next,r1494_flop_next,r1472_flop_next,b1469_flop_next,b1467_flop_next,b1465_flop_next,b1463_flop_next,b1461_flop_next,b1459_flop_next,b1457_flop_next,b1455_flop_next,b1453_flop_next,b1451_flop_next,b1449_flop_next,b1447_flop_next,b1445_flop_next,b1443_flop_next,b1441_flop_next,b1439_flop_next,r1437_flop_next,r1435_flop_next,r1433_flop_next,r1431_flop_next,r1429_flop_next,r1427_flop_next,r1425_flop_next,r1423_flop_next,r1421_flop_next,r1419_flop_next,r1417_flop_next,r1415_flop_next,r1413_flop_next,r1411_flop_next,r1409_flop_next,r1407_flop_next,b1404_flop_next,b1402_flop_next,r1400_flop_next,r1398_flop_next,r1396_flop_next,r1394_flop_next,r1388_flop_next,r1385_flop_next,b1383_flop_next,b1381_flop_next,b1379_flop_next,r1377_flop_next,r1375_flop_next,b1373_flop_next,r1365_flop_next,r1361_flop_next,r1360_flop_next,r1358_flop_next,r1336_flop_next,b1333_flop_next,b1331_flop_next,b1329_flop_next,b1327_flop_next,b1325_flop_next,b1323_flop_next,b1321_flop_next,b1319_flop_next,b1317_flop_next,b1315_flop_next,b1313_flop_next,b1311_flop_next,b1309_flop_next,b1307_flop_next,b1305_flop_next,b1303_flop_next,r1301_flop_next,r1299_flop_next,r1297_flop_next,r1295_flop_next,r1293_flop_next,r1291_flop_next,r1289_flop_next,r1287_flop_next,r1285_flop_next,r1283_flop_next,r1281_flop_next,r1279_flop_next,r1277_flop_next,r1275_flop_next,r1273_flop_next,r1271_flop_next,b1268_flop_next,b1266_flop_next,r1264_flop_next,r1262_flop_next,r1260_flop_next,r1258_flop_next,r1252_flop_next,r1249_flop_next,b1247_flop_next,b1245_flop_next,b1243_flop_next,r1241_flop_next,r1239_flop_next,b1237_flop_next,r1229_flop_next,r1225_flop_next,r1224_flop_next,r1222_flop_next,r1200_flop_next,b1197_flop_next,b1195_flop_next,b1193_flop_next,b1191_flop_next,b1189_flop_next,b1187_flop_next,b1185_flop_next,b1183_flop_next,b1181_flop_next,b1179_flop_next,b1177_flop_next,b1175_flop_next,b1173_flop_next,b1171_flop_next,b1169_flop_next,b1167_flop_next,r1165_flop_next,r1163_flop_next,r1161_flop_next,r1159_flop_next,r1157_flop_next,r1155_flop_next,r1153_flop_next,r1151_flop_next,r1149_flop_next,r1147_flop_next,r1145_flop_next,r1143_flop_next,r1141_flop_next,r1139_flop_next,r1137_flop_next,r1135_flop_next,b1132_flop_next,b1130_flop_next,r1128_flop_next,r1126_flop_next,r1124_flop_next,r1122_flop_next,r1116_flop_next,r1113_flop_next,b1111_flop_next,b1109_flop_next,b1107_flop_next,r1105_flop_next,r1103_flop_next,b1101_flop_next,r1093_flop_next,r1089_flop_next,r1088_flop_next,r1086_flop_next,r1064_flop_next,b1061_flop_next,b1059_flop_next,b1057_flop_next,b1055_flop_next,b1053_flop_next,b1051_flop_next,b1049_flop_next,b1047_flop_next,b1045_flop_next,b1043_flop_next,b1041_flop_next,b1039_flop_next,b1037_flop_next,b1035_flop_next,b1033_flop_next,b1031_flop_next,r1029_flop_next,r1027_flop_next,r1025_flop_next,r1023_flop_next,r1021_flop_next,r1019_flop_next,r1017_flop_next,r1015_flop_next,r1013_flop_next,r1011_flop_next,r1009_flop_next,r1007_flop_next,r1005_flop_next,r1003_flop_next,r1001_flop_next,r999_flop_next,b996_flop_next,b994_flop_next,r992_flop_next,r990_flop_next,r988_flop_next,r986_flop_next,r980_flop_next,r977_flop_next,b975_flop_next,b973_flop_next,b971_flop_next,r969_flop_next,r967_flop_next,b965_flop_next,r957_flop_next,r953_flop_next,r952_flop_next,r950_flop_next,r928_flop_next,b925_flop_next,b923_flop_next,b921_flop_next,b919_flop_next,b917_flop_next,b915_flop_next,b913_flop_next,b911_flop_next,b909_flop_next,b907_flop_next,b905_flop_next,b903_flop_next,b901_flop_next,b899_flop_next,b897_flop_next,b895_flop_next,r893_flop_next,r891_flop_next,r889_flop_next,r887_flop_next,r885_flop_next,r883_flop_next,r881_flop_next,r879_flop_next,r877_flop_next,r875_flop_next,r873_flop_next,r871_flop_next,r869_flop_next,r867_flop_next,r865_flop_next,r863_flop_next,b860_flop_next,b858_flop_next,r856_flop_next,r854_flop_next,r852_flop_next,r850_flop_next,r844_flop_next,r841_flop_next,b839_flop_next,b837_flop_next,b835_flop_next,r833_flop_next,r831_flop_next,b829_flop_next,r821_flop_next,r817_flop_next,r816_flop_next,r814_flop_next,r792_flop_next,b789_flop_next,b787_flop_next,b785_flop_next,b783_flop_next,b781_flop_next,b779_flop_next,b777_flop_next,b775_flop_next,b773_flop_next,b771_flop_next,b769_flop_next,b767_flop_next,b765_flop_next,b763_flop_next,b761_flop_next,b759_flop_next,r757_flop_next,r755_flop_next,r753_flop_next,r751_flop_next,r749_flop_next,r747_flop_next,r745_flop_next,r743_flop_next,r741_flop_next,r739_flop_next,r737_flop_next,r735_flop_next,r733_flop_next,r731_flop_next,r729_flop_next,r727_flop_next,b724_flop_next,b722_flop_next,r720_flop_next,r718_flop_next,r716_flop_next,r714_flop_next,r708_flop_next,r705_flop_next,b703_flop_next,b701_flop_next,b699_flop_next,r697_flop_next,r695_flop_next,b693_flop_next,r685_flop_next,r681_flop_next,r680_flop_next,r678_flop_next,r656_flop_next,b653_flop_next,b651_flop_next,b649_flop_next,b647_flop_next,b645_flop_next,b643_flop_next,b641_flop_next,b639_flop_next,b637_flop_next,b635_flop_next,b633_flop_next,b631_flop_next,b629_flop_next,b627_flop_next,b625_flop_next,b623_flop_next,r621_flop_next,r619_flop_next,r617_flop_next,r615_flop_next,r613_flop_next,r611_flop_next,r609_flop_next,r607_flop_next,r605_flop_next,r603_flop_next,r601_flop_next,r599_flop_next,r597_flop_next,r595_flop_next,r593_flop_next,r591_flop_next,b588_flop_next,b586_flop_next,r584_flop_next,r582_flop_next,r580_flop_next,r578_flop_next,r572_flop_next,r569_flop_next,r566_flop_next,b26_flop_next,b24_flop_next,b22_flop_next,r20_flop_next,r18_flop_next,b16_flop_next,r12_flop_next,r10_flop_next,r6_flop_next,r5_flop_next,r3_flop_next,statevar0_flop_next,statevar1_flop_next,statevar2_flop_next,statevar3_flop_next)
  begin
    if clk'event and clk='1' then
      input_flop <= input;
      control_flop <= control_flop_next;
      goto_L7851_flop <= goto_L7851_flop_next;
      goto_L7844_flop <= goto_L7844_flop_next;
      goto_L7806_flop <= goto_L7806_flop_next;
      goto_L7767_flop <= goto_L7767_flop_next;
      goto_L7728_flop <= goto_L7728_flop_next;
      goto_L7570_flop <= goto_L7570_flop_next;
      goto_L7690_flop <= goto_L7690_flop_next;
      goto_L7575_flop <= goto_L7575_flop_next;
      goto_L1784_flop <= goto_L1784_flop_next;
      goto_L1785_flop <= goto_L1785_flop_next;
      goto_L1638_flop <= goto_L1638_flop_next;
      goto_L1502_flop <= goto_L1502_flop_next;
      goto_L1366_flop <= goto_L1366_flop_next;
      goto_L1230_flop <= goto_L1230_flop_next;
      goto_L1094_flop <= goto_L1094_flop_next;
      goto_L958_flop <= goto_L958_flop_next;
      goto_L822_flop <= goto_L822_flop_next;
      goto_L686_flop <= goto_L686_flop_next;
      goto_L11_flop <= goto_L11_flop_next;
      goto_L13_flop <= goto_L13_flop_next;
      goto_L690_flop <= goto_L690_flop_next;
      goto_L826_flop <= goto_L826_flop_next;
      goto_L962_flop <= goto_L962_flop_next;
      goto_L1098_flop <= goto_L1098_flop_next;
      goto_L1234_flop <= goto_L1234_flop_next;
      goto_L1370_flop <= goto_L1370_flop_next;
      goto_L1506_flop <= goto_L1506_flop_next;
      goto_L1642_flop <= goto_L1642_flop_next;
      goto_L7693_flop <= goto_L7693_flop_next;
      goto_L7732_flop <= goto_L7732_flop_next;
      goto_L7771_flop <= goto_L7771_flop_next;
      goto_L7810_flop <= goto_L7810_flop_next;
      goto_L7777_flop <= goto_L7777_flop_next;
      goto_L7738_flop <= goto_L7738_flop_next;
      goto_L7699_flop <= goto_L7699_flop_next;
      goto_L1658_flop <= goto_L1658_flop_next;
      goto_L1522_flop <= goto_L1522_flop_next;
      goto_L1386_flop <= goto_L1386_flop_next;
      goto_L1250_flop <= goto_L1250_flop_next;
      goto_L1114_flop <= goto_L1114_flop_next;
      goto_L978_flop <= goto_L978_flop_next;
      goto_L842_flop <= goto_L842_flop_next;
      goto_L706_flop <= goto_L706_flop_next;
      goto_L567_flop <= goto_L567_flop_next;
      goto_L0_flop <= goto_L0_flop_next;
      goto_L7852_flop <= goto_L7852_flop_next;
      r7843_flop <= r7843_flop_next;
      r7840_flop <= r7840_flop_next;
      r7817_flop <= r7817_flop_next;
      r7814_flop <= r7814_flop_next;
      r7805_flop <= r7805_flop_next;
      r7802_flop <= r7802_flop_next;
      r7779_flop <= r7779_flop_next;
      r7776_flop <= r7776_flop_next;
      b7774_flop <= b7774_flop_next;
      r7766_flop <= r7766_flop_next;
      r7763_flop <= r7763_flop_next;
      r7740_flop <= r7740_flop_next;
      r7737_flop <= r7737_flop_next;
      b7735_flop <= b7735_flop_next;
      r7727_flop <= r7727_flop_next;
      r7724_flop <= r7724_flop_next;
      r7701_flop <= r7701_flop_next;
      r7698_flop <= r7698_flop_next;
      b7696_flop <= b7696_flop_next;
      r7679_flop <= r7679_flop_next;
      r7675_flop <= r7675_flop_next;
      r7671_flop <= r7671_flop_next;
      r7667_flop <= r7667_flop_next;
      r7663_flop <= r7663_flop_next;
      r7659_flop <= r7659_flop_next;
      r7655_flop <= r7655_flop_next;
      r7651_flop <= r7651_flop_next;
      r7647_flop <= r7647_flop_next;
      b7644_flop <= b7644_flop_next;
      b7642_flop <= b7642_flop_next;
      b7640_flop <= b7640_flop_next;
      b7638_flop <= b7638_flop_next;
      b7636_flop <= b7636_flop_next;
      b7634_flop <= b7634_flop_next;
      b7632_flop <= b7632_flop_next;
      b7630_flop <= b7630_flop_next;
      r7628_flop <= r7628_flop_next;
      r7626_flop <= r7626_flop_next;
      r7624_flop <= r7624_flop_next;
      r7622_flop <= r7622_flop_next;
      r7620_flop <= r7620_flop_next;
      r7618_flop <= r7618_flop_next;
      r7616_flop <= r7616_flop_next;
      r7614_flop <= r7614_flop_next;
      r7610_flop <= r7610_flop_next;
      b7608_flop <= b7608_flop_next;
      b7606_flop <= b7606_flop_next;
      b7604_flop <= b7604_flop_next;
      b7602_flop <= b7602_flop_next;
      b7600_flop <= b7600_flop_next;
      b7598_flop <= b7598_flop_next;
      b7596_flop <= b7596_flop_next;
      b7594_flop <= b7594_flop_next;
      r7592_flop <= r7592_flop_next;
      r7590_flop <= r7590_flop_next;
      r7588_flop <= r7588_flop_next;
      r7586_flop <= r7586_flop_next;
      r7584_flop <= r7584_flop_next;
      r7582_flop <= r7582_flop_next;
      r7580_flop <= r7580_flop_next;
      r7578_flop <= r7578_flop_next;
      r7574_flop <= r7574_flop_next;
      b7572_flop <= b7572_flop_next;
      r7569_flop <= r7569_flop_next;
      r7565_flop <= r7565_flop_next;
      r7564_flop <= r7564_flop_next;
      r7562_flop <= r7562_flop_next;
      r7558_flop <= r7558_flop_next;
      r7300_flop <= r7300_flop_next;
      r7296_flop <= r7296_flop_next;
      r7292_flop <= r7292_flop_next;
      r2874_flop <= r2874_flop_next;
      r2376_flop <= r2376_flop_next;
      r2375_flop <= r2375_flop_next;
      r2374_flop <= r2374_flop_next;
      r2371_flop <= r2371_flop_next;
      r2365_flop <= r2365_flop_next;
      r1862_flop <= r1862_flop_next;
      b1859_flop <= b1859_flop_next;
      b1857_flop <= b1857_flop_next;
      b1855_flop <= b1855_flop_next;
      b1853_flop <= b1853_flop_next;
      b1851_flop <= b1851_flop_next;
      b1849_flop <= b1849_flop_next;
      b1847_flop <= b1847_flop_next;
      b1845_flop <= b1845_flop_next;
      b1843_flop <= b1843_flop_next;
      b1841_flop <= b1841_flop_next;
      b1839_flop <= b1839_flop_next;
      b1837_flop <= b1837_flop_next;
      b1835_flop <= b1835_flop_next;
      b1833_flop <= b1833_flop_next;
      b1831_flop <= b1831_flop_next;
      b1829_flop <= b1829_flop_next;
      r1827_flop <= r1827_flop_next;
      r1825_flop <= r1825_flop_next;
      r1823_flop <= r1823_flop_next;
      r1821_flop <= r1821_flop_next;
      r1819_flop <= r1819_flop_next;
      r1817_flop <= r1817_flop_next;
      r1815_flop <= r1815_flop_next;
      r1813_flop <= r1813_flop_next;
      r1811_flop <= r1811_flop_next;
      r1809_flop <= r1809_flop_next;
      r1807_flop <= r1807_flop_next;
      r1805_flop <= r1805_flop_next;
      r1803_flop <= r1803_flop_next;
      r1801_flop <= r1801_flop_next;
      r1799_flop <= r1799_flop_next;
      r1797_flop <= r1797_flop_next;
      r1795_flop <= r1795_flop_next;
      r1792_flop <= r1792_flop_next;
      r1790_flop <= r1790_flop_next;
      r1787_flop <= r1787_flop_next;
      r1783_flop <= r1783_flop_next;
      r1779_flop <= r1779_flop_next;
      r1778_flop <= r1778_flop_next;
      r1776_flop <= r1776_flop_next;
      r1754_flop <= r1754_flop_next;
      b1751_flop <= b1751_flop_next;
      b1749_flop <= b1749_flop_next;
      b1747_flop <= b1747_flop_next;
      b1745_flop <= b1745_flop_next;
      b1743_flop <= b1743_flop_next;
      b1741_flop <= b1741_flop_next;
      b1739_flop <= b1739_flop_next;
      b1737_flop <= b1737_flop_next;
      b1735_flop <= b1735_flop_next;
      b1733_flop <= b1733_flop_next;
      b1731_flop <= b1731_flop_next;
      b1729_flop <= b1729_flop_next;
      b1727_flop <= b1727_flop_next;
      b1725_flop <= b1725_flop_next;
      b1723_flop <= b1723_flop_next;
      b1721_flop <= b1721_flop_next;
      r1719_flop <= r1719_flop_next;
      r1717_flop <= r1717_flop_next;
      r1715_flop <= r1715_flop_next;
      r1713_flop <= r1713_flop_next;
      r1711_flop <= r1711_flop_next;
      r1709_flop <= r1709_flop_next;
      r1707_flop <= r1707_flop_next;
      r1705_flop <= r1705_flop_next;
      r1703_flop <= r1703_flop_next;
      r1701_flop <= r1701_flop_next;
      r1699_flop <= r1699_flop_next;
      r1697_flop <= r1697_flop_next;
      r1695_flop <= r1695_flop_next;
      r1693_flop <= r1693_flop_next;
      r1691_flop <= r1691_flop_next;
      r1689_flop <= r1689_flop_next;
      b1686_flop <= b1686_flop_next;
      b1684_flop <= b1684_flop_next;
      r1682_flop <= r1682_flop_next;
      r1680_flop <= r1680_flop_next;
      r1678_flop <= r1678_flop_next;
      r1676_flop <= r1676_flop_next;
      r1670_flop <= r1670_flop_next;
      r1667_flop <= r1667_flop_next;
      r1663_flop <= r1663_flop_next;
      r1659_flop <= r1659_flop_next;
      r1657_flop <= r1657_flop_next;
      b1655_flop <= b1655_flop_next;
      b1653_flop <= b1653_flop_next;
      b1651_flop <= b1651_flop_next;
      r1649_flop <= r1649_flop_next;
      r1647_flop <= r1647_flop_next;
      b1645_flop <= b1645_flop_next;
      r1637_flop <= r1637_flop_next;
      r1633_flop <= r1633_flop_next;
      r1632_flop <= r1632_flop_next;
      r1630_flop <= r1630_flop_next;
      r1608_flop <= r1608_flop_next;
      b1605_flop <= b1605_flop_next;
      b1603_flop <= b1603_flop_next;
      b1601_flop <= b1601_flop_next;
      b1599_flop <= b1599_flop_next;
      b1597_flop <= b1597_flop_next;
      b1595_flop <= b1595_flop_next;
      b1593_flop <= b1593_flop_next;
      b1591_flop <= b1591_flop_next;
      b1589_flop <= b1589_flop_next;
      b1587_flop <= b1587_flop_next;
      b1585_flop <= b1585_flop_next;
      b1583_flop <= b1583_flop_next;
      b1581_flop <= b1581_flop_next;
      b1579_flop <= b1579_flop_next;
      b1577_flop <= b1577_flop_next;
      b1575_flop <= b1575_flop_next;
      r1573_flop <= r1573_flop_next;
      r1571_flop <= r1571_flop_next;
      r1569_flop <= r1569_flop_next;
      r1567_flop <= r1567_flop_next;
      r1565_flop <= r1565_flop_next;
      r1563_flop <= r1563_flop_next;
      r1561_flop <= r1561_flop_next;
      r1559_flop <= r1559_flop_next;
      r1557_flop <= r1557_flop_next;
      r1555_flop <= r1555_flop_next;
      r1553_flop <= r1553_flop_next;
      r1551_flop <= r1551_flop_next;
      r1549_flop <= r1549_flop_next;
      r1547_flop <= r1547_flop_next;
      r1545_flop <= r1545_flop_next;
      r1543_flop <= r1543_flop_next;
      b1540_flop <= b1540_flop_next;
      b1538_flop <= b1538_flop_next;
      r1536_flop <= r1536_flop_next;
      r1534_flop <= r1534_flop_next;
      r1532_flop <= r1532_flop_next;
      r1530_flop <= r1530_flop_next;
      r1524_flop <= r1524_flop_next;
      r1521_flop <= r1521_flop_next;
      b1519_flop <= b1519_flop_next;
      b1517_flop <= b1517_flop_next;
      b1515_flop <= b1515_flop_next;
      r1513_flop <= r1513_flop_next;
      r1511_flop <= r1511_flop_next;
      b1509_flop <= b1509_flop_next;
      r1501_flop <= r1501_flop_next;
      r1497_flop <= r1497_flop_next;
      r1496_flop <= r1496_flop_next;
      r1494_flop <= r1494_flop_next;
      r1472_flop <= r1472_flop_next;
      b1469_flop <= b1469_flop_next;
      b1467_flop <= b1467_flop_next;
      b1465_flop <= b1465_flop_next;
      b1463_flop <= b1463_flop_next;
      b1461_flop <= b1461_flop_next;
      b1459_flop <= b1459_flop_next;
      b1457_flop <= b1457_flop_next;
      b1455_flop <= b1455_flop_next;
      b1453_flop <= b1453_flop_next;
      b1451_flop <= b1451_flop_next;
      b1449_flop <= b1449_flop_next;
      b1447_flop <= b1447_flop_next;
      b1445_flop <= b1445_flop_next;
      b1443_flop <= b1443_flop_next;
      b1441_flop <= b1441_flop_next;
      b1439_flop <= b1439_flop_next;
      r1437_flop <= r1437_flop_next;
      r1435_flop <= r1435_flop_next;
      r1433_flop <= r1433_flop_next;
      r1431_flop <= r1431_flop_next;
      r1429_flop <= r1429_flop_next;
      r1427_flop <= r1427_flop_next;
      r1425_flop <= r1425_flop_next;
      r1423_flop <= r1423_flop_next;
      r1421_flop <= r1421_flop_next;
      r1419_flop <= r1419_flop_next;
      r1417_flop <= r1417_flop_next;
      r1415_flop <= r1415_flop_next;
      r1413_flop <= r1413_flop_next;
      r1411_flop <= r1411_flop_next;
      r1409_flop <= r1409_flop_next;
      r1407_flop <= r1407_flop_next;
      b1404_flop <= b1404_flop_next;
      b1402_flop <= b1402_flop_next;
      r1400_flop <= r1400_flop_next;
      r1398_flop <= r1398_flop_next;
      r1396_flop <= r1396_flop_next;
      r1394_flop <= r1394_flop_next;
      r1388_flop <= r1388_flop_next;
      r1385_flop <= r1385_flop_next;
      b1383_flop <= b1383_flop_next;
      b1381_flop <= b1381_flop_next;
      b1379_flop <= b1379_flop_next;
      r1377_flop <= r1377_flop_next;
      r1375_flop <= r1375_flop_next;
      b1373_flop <= b1373_flop_next;
      r1365_flop <= r1365_flop_next;
      r1361_flop <= r1361_flop_next;
      r1360_flop <= r1360_flop_next;
      r1358_flop <= r1358_flop_next;
      r1336_flop <= r1336_flop_next;
      b1333_flop <= b1333_flop_next;
      b1331_flop <= b1331_flop_next;
      b1329_flop <= b1329_flop_next;
      b1327_flop <= b1327_flop_next;
      b1325_flop <= b1325_flop_next;
      b1323_flop <= b1323_flop_next;
      b1321_flop <= b1321_flop_next;
      b1319_flop <= b1319_flop_next;
      b1317_flop <= b1317_flop_next;
      b1315_flop <= b1315_flop_next;
      b1313_flop <= b1313_flop_next;
      b1311_flop <= b1311_flop_next;
      b1309_flop <= b1309_flop_next;
      b1307_flop <= b1307_flop_next;
      b1305_flop <= b1305_flop_next;
      b1303_flop <= b1303_flop_next;
      r1301_flop <= r1301_flop_next;
      r1299_flop <= r1299_flop_next;
      r1297_flop <= r1297_flop_next;
      r1295_flop <= r1295_flop_next;
      r1293_flop <= r1293_flop_next;
      r1291_flop <= r1291_flop_next;
      r1289_flop <= r1289_flop_next;
      r1287_flop <= r1287_flop_next;
      r1285_flop <= r1285_flop_next;
      r1283_flop <= r1283_flop_next;
      r1281_flop <= r1281_flop_next;
      r1279_flop <= r1279_flop_next;
      r1277_flop <= r1277_flop_next;
      r1275_flop <= r1275_flop_next;
      r1273_flop <= r1273_flop_next;
      r1271_flop <= r1271_flop_next;
      b1268_flop <= b1268_flop_next;
      b1266_flop <= b1266_flop_next;
      r1264_flop <= r1264_flop_next;
      r1262_flop <= r1262_flop_next;
      r1260_flop <= r1260_flop_next;
      r1258_flop <= r1258_flop_next;
      r1252_flop <= r1252_flop_next;
      r1249_flop <= r1249_flop_next;
      b1247_flop <= b1247_flop_next;
      b1245_flop <= b1245_flop_next;
      b1243_flop <= b1243_flop_next;
      r1241_flop <= r1241_flop_next;
      r1239_flop <= r1239_flop_next;
      b1237_flop <= b1237_flop_next;
      r1229_flop <= r1229_flop_next;
      r1225_flop <= r1225_flop_next;
      r1224_flop <= r1224_flop_next;
      r1222_flop <= r1222_flop_next;
      r1200_flop <= r1200_flop_next;
      b1197_flop <= b1197_flop_next;
      b1195_flop <= b1195_flop_next;
      b1193_flop <= b1193_flop_next;
      b1191_flop <= b1191_flop_next;
      b1189_flop <= b1189_flop_next;
      b1187_flop <= b1187_flop_next;
      b1185_flop <= b1185_flop_next;
      b1183_flop <= b1183_flop_next;
      b1181_flop <= b1181_flop_next;
      b1179_flop <= b1179_flop_next;
      b1177_flop <= b1177_flop_next;
      b1175_flop <= b1175_flop_next;
      b1173_flop <= b1173_flop_next;
      b1171_flop <= b1171_flop_next;
      b1169_flop <= b1169_flop_next;
      b1167_flop <= b1167_flop_next;
      r1165_flop <= r1165_flop_next;
      r1163_flop <= r1163_flop_next;
      r1161_flop <= r1161_flop_next;
      r1159_flop <= r1159_flop_next;
      r1157_flop <= r1157_flop_next;
      r1155_flop <= r1155_flop_next;
      r1153_flop <= r1153_flop_next;
      r1151_flop <= r1151_flop_next;
      r1149_flop <= r1149_flop_next;
      r1147_flop <= r1147_flop_next;
      r1145_flop <= r1145_flop_next;
      r1143_flop <= r1143_flop_next;
      r1141_flop <= r1141_flop_next;
      r1139_flop <= r1139_flop_next;
      r1137_flop <= r1137_flop_next;
      r1135_flop <= r1135_flop_next;
      b1132_flop <= b1132_flop_next;
      b1130_flop <= b1130_flop_next;
      r1128_flop <= r1128_flop_next;
      r1126_flop <= r1126_flop_next;
      r1124_flop <= r1124_flop_next;
      r1122_flop <= r1122_flop_next;
      r1116_flop <= r1116_flop_next;
      r1113_flop <= r1113_flop_next;
      b1111_flop <= b1111_flop_next;
      b1109_flop <= b1109_flop_next;
      b1107_flop <= b1107_flop_next;
      r1105_flop <= r1105_flop_next;
      r1103_flop <= r1103_flop_next;
      b1101_flop <= b1101_flop_next;
      r1093_flop <= r1093_flop_next;
      r1089_flop <= r1089_flop_next;
      r1088_flop <= r1088_flop_next;
      r1086_flop <= r1086_flop_next;
      r1064_flop <= r1064_flop_next;
      b1061_flop <= b1061_flop_next;
      b1059_flop <= b1059_flop_next;
      b1057_flop <= b1057_flop_next;
      b1055_flop <= b1055_flop_next;
      b1053_flop <= b1053_flop_next;
      b1051_flop <= b1051_flop_next;
      b1049_flop <= b1049_flop_next;
      b1047_flop <= b1047_flop_next;
      b1045_flop <= b1045_flop_next;
      b1043_flop <= b1043_flop_next;
      b1041_flop <= b1041_flop_next;
      b1039_flop <= b1039_flop_next;
      b1037_flop <= b1037_flop_next;
      b1035_flop <= b1035_flop_next;
      b1033_flop <= b1033_flop_next;
      b1031_flop <= b1031_flop_next;
      r1029_flop <= r1029_flop_next;
      r1027_flop <= r1027_flop_next;
      r1025_flop <= r1025_flop_next;
      r1023_flop <= r1023_flop_next;
      r1021_flop <= r1021_flop_next;
      r1019_flop <= r1019_flop_next;
      r1017_flop <= r1017_flop_next;
      r1015_flop <= r1015_flop_next;
      r1013_flop <= r1013_flop_next;
      r1011_flop <= r1011_flop_next;
      r1009_flop <= r1009_flop_next;
      r1007_flop <= r1007_flop_next;
      r1005_flop <= r1005_flop_next;
      r1003_flop <= r1003_flop_next;
      r1001_flop <= r1001_flop_next;
      r999_flop <= r999_flop_next;
      b996_flop <= b996_flop_next;
      b994_flop <= b994_flop_next;
      r992_flop <= r992_flop_next;
      r990_flop <= r990_flop_next;
      r988_flop <= r988_flop_next;
      r986_flop <= r986_flop_next;
      r980_flop <= r980_flop_next;
      r977_flop <= r977_flop_next;
      b975_flop <= b975_flop_next;
      b973_flop <= b973_flop_next;
      b971_flop <= b971_flop_next;
      r969_flop <= r969_flop_next;
      r967_flop <= r967_flop_next;
      b965_flop <= b965_flop_next;
      r957_flop <= r957_flop_next;
      r953_flop <= r953_flop_next;
      r952_flop <= r952_flop_next;
      r950_flop <= r950_flop_next;
      r928_flop <= r928_flop_next;
      b925_flop <= b925_flop_next;
      b923_flop <= b923_flop_next;
      b921_flop <= b921_flop_next;
      b919_flop <= b919_flop_next;
      b917_flop <= b917_flop_next;
      b915_flop <= b915_flop_next;
      b913_flop <= b913_flop_next;
      b911_flop <= b911_flop_next;
      b909_flop <= b909_flop_next;
      b907_flop <= b907_flop_next;
      b905_flop <= b905_flop_next;
      b903_flop <= b903_flop_next;
      b901_flop <= b901_flop_next;
      b899_flop <= b899_flop_next;
      b897_flop <= b897_flop_next;
      b895_flop <= b895_flop_next;
      r893_flop <= r893_flop_next;
      r891_flop <= r891_flop_next;
      r889_flop <= r889_flop_next;
      r887_flop <= r887_flop_next;
      r885_flop <= r885_flop_next;
      r883_flop <= r883_flop_next;
      r881_flop <= r881_flop_next;
      r879_flop <= r879_flop_next;
      r877_flop <= r877_flop_next;
      r875_flop <= r875_flop_next;
      r873_flop <= r873_flop_next;
      r871_flop <= r871_flop_next;
      r869_flop <= r869_flop_next;
      r867_flop <= r867_flop_next;
      r865_flop <= r865_flop_next;
      r863_flop <= r863_flop_next;
      b860_flop <= b860_flop_next;
      b858_flop <= b858_flop_next;
      r856_flop <= r856_flop_next;
      r854_flop <= r854_flop_next;
      r852_flop <= r852_flop_next;
      r850_flop <= r850_flop_next;
      r844_flop <= r844_flop_next;
      r841_flop <= r841_flop_next;
      b839_flop <= b839_flop_next;
      b837_flop <= b837_flop_next;
      b835_flop <= b835_flop_next;
      r833_flop <= r833_flop_next;
      r831_flop <= r831_flop_next;
      b829_flop <= b829_flop_next;
      r821_flop <= r821_flop_next;
      r817_flop <= r817_flop_next;
      r816_flop <= r816_flop_next;
      r814_flop <= r814_flop_next;
      r792_flop <= r792_flop_next;
      b789_flop <= b789_flop_next;
      b787_flop <= b787_flop_next;
      b785_flop <= b785_flop_next;
      b783_flop <= b783_flop_next;
      b781_flop <= b781_flop_next;
      b779_flop <= b779_flop_next;
      b777_flop <= b777_flop_next;
      b775_flop <= b775_flop_next;
      b773_flop <= b773_flop_next;
      b771_flop <= b771_flop_next;
      b769_flop <= b769_flop_next;
      b767_flop <= b767_flop_next;
      b765_flop <= b765_flop_next;
      b763_flop <= b763_flop_next;
      b761_flop <= b761_flop_next;
      b759_flop <= b759_flop_next;
      r757_flop <= r757_flop_next;
      r755_flop <= r755_flop_next;
      r753_flop <= r753_flop_next;
      r751_flop <= r751_flop_next;
      r749_flop <= r749_flop_next;
      r747_flop <= r747_flop_next;
      r745_flop <= r745_flop_next;
      r743_flop <= r743_flop_next;
      r741_flop <= r741_flop_next;
      r739_flop <= r739_flop_next;
      r737_flop <= r737_flop_next;
      r735_flop <= r735_flop_next;
      r733_flop <= r733_flop_next;
      r731_flop <= r731_flop_next;
      r729_flop <= r729_flop_next;
      r727_flop <= r727_flop_next;
      b724_flop <= b724_flop_next;
      b722_flop <= b722_flop_next;
      r720_flop <= r720_flop_next;
      r718_flop <= r718_flop_next;
      r716_flop <= r716_flop_next;
      r714_flop <= r714_flop_next;
      r708_flop <= r708_flop_next;
      r705_flop <= r705_flop_next;
      b703_flop <= b703_flop_next;
      b701_flop <= b701_flop_next;
      b699_flop <= b699_flop_next;
      r697_flop <= r697_flop_next;
      r695_flop <= r695_flop_next;
      b693_flop <= b693_flop_next;
      r685_flop <= r685_flop_next;
      r681_flop <= r681_flop_next;
      r680_flop <= r680_flop_next;
      r678_flop <= r678_flop_next;
      r656_flop <= r656_flop_next;
      b653_flop <= b653_flop_next;
      b651_flop <= b651_flop_next;
      b649_flop <= b649_flop_next;
      b647_flop <= b647_flop_next;
      b645_flop <= b645_flop_next;
      b643_flop <= b643_flop_next;
      b641_flop <= b641_flop_next;
      b639_flop <= b639_flop_next;
      b637_flop <= b637_flop_next;
      b635_flop <= b635_flop_next;
      b633_flop <= b633_flop_next;
      b631_flop <= b631_flop_next;
      b629_flop <= b629_flop_next;
      b627_flop <= b627_flop_next;
      b625_flop <= b625_flop_next;
      b623_flop <= b623_flop_next;
      r621_flop <= r621_flop_next;
      r619_flop <= r619_flop_next;
      r617_flop <= r617_flop_next;
      r615_flop <= r615_flop_next;
      r613_flop <= r613_flop_next;
      r611_flop <= r611_flop_next;
      r609_flop <= r609_flop_next;
      r607_flop <= r607_flop_next;
      r605_flop <= r605_flop_next;
      r603_flop <= r603_flop_next;
      r601_flop <= r601_flop_next;
      r599_flop <= r599_flop_next;
      r597_flop <= r597_flop_next;
      r595_flop <= r595_flop_next;
      r593_flop <= r593_flop_next;
      r591_flop <= r591_flop_next;
      b588_flop <= b588_flop_next;
      b586_flop <= b586_flop_next;
      r584_flop <= r584_flop_next;
      r582_flop <= r582_flop_next;
      r580_flop <= r580_flop_next;
      r578_flop <= r578_flop_next;
      r572_flop <= r572_flop_next;
      r569_flop <= r569_flop_next;
      r566_flop <= r566_flop_next;
      b26_flop <= b26_flop_next;
      b24_flop <= b24_flop_next;
      b22_flop <= b22_flop_next;
      r20_flop <= r20_flop_next;
      r18_flop <= r18_flop_next;
      b16_flop <= b16_flop_next;
      r12_flop <= r12_flop_next;
      r10_flop <= r10_flop_next;
      r6_flop <= r6_flop_next;
      r5_flop <= r5_flop_next;
      r3_flop <= r3_flop_next;
      statevar0_flop <= statevar0_flop_next;
      statevar1_flop <= statevar1_flop_next;
      statevar2_flop <= statevar2_flop_next;
      statevar3_flop <= statevar3_flop_next;
    end if;
  end process;

end behavioral;
