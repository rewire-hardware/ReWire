library ieee;
use ieee.std_logic_1164.all;
-- Comment out the following line if VHDL primitives are not in use.
use work.prims.all;
entity rewire is
  Port ( clk : in std_logic ;
         input : in std_logic_vector (0 to 513);
         output : out std_logic_vector (0 to 257));
end rewire;

architecture behavioral of rewire is
  type control_state is (STATE0,STATE11,STATE585,STATE6110,STATE6264,STATE6280);
  function rewire_Main.seed_1671(r1672 : std_logic_vector) return std_logic_vector;
  function rewire_MetaprogrammingRW.wc67178f2_6022 return std_logic_vector;
  function rewire_MetaprogrammingRW.wbef9a3f7_5953 return std_logic_vector;
  function rewire_MetaprogrammingRW.wa4506ceb_5884 return std_logic_vector;
  function rewire_MetaprogrammingRW.w90befffa_5815 return std_logic_vector;
  function rewire_MetaprogrammingRW.w8cc70208_5746 return std_logic_vector;
  function rewire_MetaprogrammingRW.w84c87814_5677 return std_logic_vector;
  function rewire_MetaprogrammingRW.w78a5636f_5608 return std_logic_vector;
  function rewire_MetaprogrammingRW.w748f82ee_5539 return std_logic_vector;
  function rewire_MetaprogrammingRW.w682e6ff3_5470 return std_logic_vector;
  function rewire_MetaprogrammingRW.w5b9cca4f_5401 return std_logic_vector;
  function rewire_MetaprogrammingRW.w4ed8aa4a_5332 return std_logic_vector;
  function rewire_MetaprogrammingRW.w391c0cb3_5263 return std_logic_vector;
  function rewire_MetaprogrammingRW.w34b0bcb5_5194 return std_logic_vector;
  function rewire_MetaprogrammingRW.w2748774c_5125 return std_logic_vector;
  function rewire_MetaprogrammingRW.w1e376c08_5056 return std_logic_vector;
  function rewire_MetaprogrammingRW.w19a4c116_4987 return std_logic_vector;
  function rewire_MetaprogrammingRW.w106aa070_4918 return std_logic_vector;
  function rewire_MetaprogrammingRW.wf40e3585_4849 return std_logic_vector;
  function rewire_MetaprogrammingRW.wd6990624_4780 return std_logic_vector;
  function rewire_MetaprogrammingRW.wd192e819_4711 return std_logic_vector;
  function rewire_MetaprogrammingRW.wc76c51a3_4642 return std_logic_vector;
  function rewire_MetaprogrammingRW.wc24b8b70_4573 return std_logic_vector;
  function rewire_MetaprogrammingRW.wa81a664b_4504 return std_logic_vector;
  function rewire_MetaprogrammingRW.wa2bfe8a1_4435 return std_logic_vector;
  function rewire_MetaprogrammingRW.w92722c85_4366 return std_logic_vector;
  function rewire_MetaprogrammingRW.w81c2c92e_4297 return std_logic_vector;
  function rewire_MetaprogrammingRW.w766a0abb_4228 return std_logic_vector;
  function rewire_MetaprogrammingRW.w650a7354_4159 return std_logic_vector;
  function rewire_MetaprogrammingRW.w53380d13_4090 return std_logic_vector;
  function rewire_MetaprogrammingRW.w4d2c6dfc_4021 return std_logic_vector;
  function rewire_MetaprogrammingRW.w2e1b2138_3952 return std_logic_vector;
  function rewire_MetaprogrammingRW.w27b70a85_3883 return std_logic_vector;
  function rewire_MetaprogrammingRW.w14292967_3814 return std_logic_vector;
  function rewire_MetaprogrammingRW.w06ca6351_3745 return std_logic_vector;
  function rewire_MetaprogrammingRW.wd5a79147_3676 return std_logic_vector;
  function rewire_MetaprogrammingRW.wc6e00bf3_3607 return std_logic_vector;
  function rewire_MetaprogrammingRW.wbf597fc7_3538 return std_logic_vector;
  function rewire_MetaprogrammingRW.wb00327c8_3469 return std_logic_vector;
  function rewire_MetaprogrammingRW.wa831c66d_3400 return std_logic_vector;
  function rewire_MetaprogrammingRW.w983e5152_3331 return std_logic_vector;
  function rewire_MetaprogrammingRW.w76f988da_3262 return std_logic_vector;
  function rewire_MetaprogrammingRW.w5cb0a9dc_3193 return std_logic_vector;
  function rewire_MetaprogrammingRW.w4a7484aa_3124 return std_logic_vector;
  function rewire_MetaprogrammingRW.w2de92c6f_3055 return std_logic_vector;
  function rewire_MetaprogrammingRW.w240ca1cc_2986 return std_logic_vector;
  function rewire_MetaprogrammingRW.w0fc19dc6_2917 return std_logic_vector;
  function rewire_MetaprogrammingRW.wefbe4786_2848 return std_logic_vector;
  function rewire_MetaprogrammingRW.we49b69c1_2779 return std_logic_vector;
  function rewire_MetaprogrammingRW.wc19bf174_2710 return std_logic_vector;
  function rewire_MetaprogrammingRW.w9bdc06a7_2641 return std_logic_vector;
  function rewire_MetaprogrammingRW.w80deb1fe_2572 return std_logic_vector;
  function rewire_MetaprogrammingRW.w72be5d74_2503 return std_logic_vector;
  function rewire_MetaprogrammingRW.w550c7dc3_2434 return std_logic_vector;
  function rewire_MetaprogrammingRW.w243185be_2365 return std_logic_vector;
  function rewire_MetaprogrammingRW.w12835b01_2296 return std_logic_vector;
  function rewire_MetaprogrammingRW.wd807aa98_2227 return std_logic_vector;
  function rewire_MetaprogrammingRW.wab1c5ed5_2158 return std_logic_vector;
  function rewire_MetaprogrammingRW.w923f82a4_2089 return std_logic_vector;
  function rewire_MetaprogrammingRW.w59f111f1_2020 return std_logic_vector;
  function rewire_MetaprogrammingRW.w3956c25b_1951 return std_logic_vector;
  function rewire_MetaprogrammingRW.we9b5dba5_1882 return std_logic_vector;
  function rewire_MetaprogrammingRW.wb5c0fbcf_1813 return std_logic_vector;
  function rewire_MetaprogrammingRW.w71374491_1744 return std_logic_vector;
  function rewire_MetaprogrammingRW.w428a2f98_1675 return std_logic_vector;
  function rewire_Main.step256_1171(r1172 : std_logic_vector ; r1173 : std_logic_vector ; r1174 : std_logic_vector) return std_logic_vector;
  function rewire_Main.maj_1652(r1653 : std_logic_vector ; r1654 : std_logic_vector ; r1655 : std_logic_vector) return std_logic_vector;
  function rewire_Main.bigsigma0_1434(r1435 : std_logic_vector) return std_logic_vector;
  function rewire_RWPrelude.rotateR22_1579(r1580 : std_logic_vector) return std_logic_vector;
  function rewire_RWPrelude.rotateR13_1507(r1508 : std_logic_vector) return std_logic_vector;
  function rewire_RWPrelude.rotateR2_1436(r1437 : std_logic_vector) return std_logic_vector;
  function rewire_Main.ch_1421(r1422 : std_logic_vector ; r1423 : std_logic_vector ; r1424 : std_logic_vector) return std_logic_vector;
  function rewire_Main.bigsigma1_1203(r1204 : std_logic_vector) return std_logic_vector;
  function rewire_RWPrelude.rotateR25_1348(r1349 : std_logic_vector) return std_logic_vector;
  function rewire_RWPrelude.rotateR11_1276(r1277 : std_logic_vector) return std_logic_vector;
  function rewire_RWPrelude.rotateR6_1205(r1206 : std_logic_vector) return std_logic_vector;
  function rewire_Main.updateSched_659(r660 : std_logic_vector) return std_logic_vector;
  function rewire_Main.sigma0_936(r937 : std_logic_vector) return std_logic_vector;
  function rewire_RWPrelude.shiftR3_1081(r1082 : std_logic_vector) return std_logic_vector;
  function rewire_RWPrelude.rotateR18_1009(r1010 : std_logic_vector) return std_logic_vector;
  function rewire_RWPrelude.rotateR7_938(r939 : std_logic_vector) return std_logic_vector;
  function rewire_Main.sigma1_697(r698 : std_logic_vector) return std_logic_vector;
  function rewire_RWPrelude.shiftR10_842(r843 : std_logic_vector) return std_logic_vector;
  function rewire_RWPrelude.rotateR19_770(r771 : std_logic_vector) return std_logic_vector;
  function rewire_RWPrelude.rotateR17_699(r700 : std_logic_vector) return std_logic_vector;
  function rewire_Main.initialSHA256State_24 return std_logic_vector;
  function rewire_MetaprogrammingRW.w5be0cd19_495 return std_logic_vector;
  function rewire_MetaprogrammingRW.w1f83d9ab_428 return std_logic_vector;
  function rewire_MetaprogrammingRW.w9b05688c_361 return std_logic_vector;
  function rewire_MetaprogrammingRW.w510e527f_294 return std_logic_vector;
  function rewire_MetaprogrammingRW.wa54ff53a_227 return std_logic_vector;
  function rewire_MetaprogrammingRW.w3c6ef372_160 return std_logic_vector;
  function rewire_MetaprogrammingRW.wbb67ae85_93 return std_logic_vector;
  function rewire_MetaprogrammingRW.w6a09e667_26 return std_logic_vector;
  function rewire_Main.seed_1671(r1672 : std_logic_vector) return std_logic_vector
  is
    variable r6088 : std_logic_vector(0 to 31) := (others => '0');
    variable b6021 : boolean := false;
    variable r6020 : std_logic_vector(0 to 31) := (others => '0');
    variable r6019 : std_logic_vector(0 to 31) := (others => '0');
    variable b5952 : boolean := false;
    variable r5951 : std_logic_vector(0 to 31) := (others => '0');
    variable r5950 : std_logic_vector(0 to 31) := (others => '0');
    variable b5883 : boolean := false;
    variable r5882 : std_logic_vector(0 to 31) := (others => '0');
    variable r5881 : std_logic_vector(0 to 31) := (others => '0');
    variable b5814 : boolean := false;
    variable r5813 : std_logic_vector(0 to 31) := (others => '0');
    variable r5812 : std_logic_vector(0 to 31) := (others => '0');
    variable b5745 : boolean := false;
    variable r5744 : std_logic_vector(0 to 31) := (others => '0');
    variable r5743 : std_logic_vector(0 to 31) := (others => '0');
    variable b5676 : boolean := false;
    variable r5675 : std_logic_vector(0 to 31) := (others => '0');
    variable r5674 : std_logic_vector(0 to 31) := (others => '0');
    variable b5607 : boolean := false;
    variable r5606 : std_logic_vector(0 to 31) := (others => '0');
    variable r5605 : std_logic_vector(0 to 31) := (others => '0');
    variable b5538 : boolean := false;
    variable r5537 : std_logic_vector(0 to 31) := (others => '0');
    variable r5536 : std_logic_vector(0 to 31) := (others => '0');
    variable b5469 : boolean := false;
    variable r5468 : std_logic_vector(0 to 31) := (others => '0');
    variable r5467 : std_logic_vector(0 to 31) := (others => '0');
    variable b5400 : boolean := false;
    variable r5399 : std_logic_vector(0 to 31) := (others => '0');
    variable r5398 : std_logic_vector(0 to 31) := (others => '0');
    variable b5331 : boolean := false;
    variable r5330 : std_logic_vector(0 to 31) := (others => '0');
    variable r5329 : std_logic_vector(0 to 31) := (others => '0');
    variable b5262 : boolean := false;
    variable r5261 : std_logic_vector(0 to 31) := (others => '0');
    variable r5260 : std_logic_vector(0 to 31) := (others => '0');
    variable b5193 : boolean := false;
    variable r5192 : std_logic_vector(0 to 31) := (others => '0');
    variable r5191 : std_logic_vector(0 to 31) := (others => '0');
    variable b5124 : boolean := false;
    variable r5123 : std_logic_vector(0 to 31) := (others => '0');
    variable r5122 : std_logic_vector(0 to 31) := (others => '0');
    variable b5055 : boolean := false;
    variable r5054 : std_logic_vector(0 to 31) := (others => '0');
    variable r5053 : std_logic_vector(0 to 31) := (others => '0');
    variable b4986 : boolean := false;
    variable r4985 : std_logic_vector(0 to 31) := (others => '0');
    variable r4984 : std_logic_vector(0 to 31) := (others => '0');
    variable b4917 : boolean := false;
    variable r4916 : std_logic_vector(0 to 31) := (others => '0');
    variable r4915 : std_logic_vector(0 to 31) := (others => '0');
    variable b4848 : boolean := false;
    variable r4847 : std_logic_vector(0 to 31) := (others => '0');
    variable r4846 : std_logic_vector(0 to 31) := (others => '0');
    variable b4779 : boolean := false;
    variable r4778 : std_logic_vector(0 to 31) := (others => '0');
    variable r4777 : std_logic_vector(0 to 31) := (others => '0');
    variable b4710 : boolean := false;
    variable r4709 : std_logic_vector(0 to 31) := (others => '0');
    variable r4708 : std_logic_vector(0 to 31) := (others => '0');
    variable b4641 : boolean := false;
    variable r4640 : std_logic_vector(0 to 31) := (others => '0');
    variable r4639 : std_logic_vector(0 to 31) := (others => '0');
    variable b4572 : boolean := false;
    variable r4571 : std_logic_vector(0 to 31) := (others => '0');
    variable r4570 : std_logic_vector(0 to 31) := (others => '0');
    variable b4503 : boolean := false;
    variable r4502 : std_logic_vector(0 to 31) := (others => '0');
    variable r4501 : std_logic_vector(0 to 31) := (others => '0');
    variable b4434 : boolean := false;
    variable r4433 : std_logic_vector(0 to 31) := (others => '0');
    variable r4432 : std_logic_vector(0 to 31) := (others => '0');
    variable b4365 : boolean := false;
    variable r4364 : std_logic_vector(0 to 31) := (others => '0');
    variable r4363 : std_logic_vector(0 to 31) := (others => '0');
    variable b4296 : boolean := false;
    variable r4295 : std_logic_vector(0 to 31) := (others => '0');
    variable r4294 : std_logic_vector(0 to 31) := (others => '0');
    variable b4227 : boolean := false;
    variable r4226 : std_logic_vector(0 to 31) := (others => '0');
    variable r4225 : std_logic_vector(0 to 31) := (others => '0');
    variable b4158 : boolean := false;
    variable r4157 : std_logic_vector(0 to 31) := (others => '0');
    variable r4156 : std_logic_vector(0 to 31) := (others => '0');
    variable b4089 : boolean := false;
    variable r4088 : std_logic_vector(0 to 31) := (others => '0');
    variable r4087 : std_logic_vector(0 to 31) := (others => '0');
    variable b4020 : boolean := false;
    variable r4019 : std_logic_vector(0 to 31) := (others => '0');
    variable r4018 : std_logic_vector(0 to 31) := (others => '0');
    variable b3951 : boolean := false;
    variable r3950 : std_logic_vector(0 to 31) := (others => '0');
    variable r3949 : std_logic_vector(0 to 31) := (others => '0');
    variable b3882 : boolean := false;
    variable r3881 : std_logic_vector(0 to 31) := (others => '0');
    variable r3880 : std_logic_vector(0 to 31) := (others => '0');
    variable b3813 : boolean := false;
    variable r3812 : std_logic_vector(0 to 31) := (others => '0');
    variable r3811 : std_logic_vector(0 to 31) := (others => '0');
    variable b3744 : boolean := false;
    variable r3743 : std_logic_vector(0 to 31) := (others => '0');
    variable r3742 : std_logic_vector(0 to 31) := (others => '0');
    variable b3675 : boolean := false;
    variable r3674 : std_logic_vector(0 to 31) := (others => '0');
    variable r3673 : std_logic_vector(0 to 31) := (others => '0');
    variable b3606 : boolean := false;
    variable r3605 : std_logic_vector(0 to 31) := (others => '0');
    variable r3604 : std_logic_vector(0 to 31) := (others => '0');
    variable b3537 : boolean := false;
    variable r3536 : std_logic_vector(0 to 31) := (others => '0');
    variable r3535 : std_logic_vector(0 to 31) := (others => '0');
    variable b3468 : boolean := false;
    variable r3467 : std_logic_vector(0 to 31) := (others => '0');
    variable r3466 : std_logic_vector(0 to 31) := (others => '0');
    variable b3399 : boolean := false;
    variable r3398 : std_logic_vector(0 to 31) := (others => '0');
    variable r3397 : std_logic_vector(0 to 31) := (others => '0');
    variable b3330 : boolean := false;
    variable r3329 : std_logic_vector(0 to 31) := (others => '0');
    variable r3328 : std_logic_vector(0 to 31) := (others => '0');
    variable b3261 : boolean := false;
    variable r3260 : std_logic_vector(0 to 31) := (others => '0');
    variable r3259 : std_logic_vector(0 to 31) := (others => '0');
    variable b3192 : boolean := false;
    variable r3191 : std_logic_vector(0 to 31) := (others => '0');
    variable r3190 : std_logic_vector(0 to 31) := (others => '0');
    variable b3123 : boolean := false;
    variable r3122 : std_logic_vector(0 to 31) := (others => '0');
    variable r3121 : std_logic_vector(0 to 31) := (others => '0');
    variable b3054 : boolean := false;
    variable r3053 : std_logic_vector(0 to 31) := (others => '0');
    variable r3052 : std_logic_vector(0 to 31) := (others => '0');
    variable b2985 : boolean := false;
    variable r2984 : std_logic_vector(0 to 31) := (others => '0');
    variable r2983 : std_logic_vector(0 to 31) := (others => '0');
    variable b2916 : boolean := false;
    variable r2915 : std_logic_vector(0 to 31) := (others => '0');
    variable r2914 : std_logic_vector(0 to 31) := (others => '0');
    variable b2847 : boolean := false;
    variable r2846 : std_logic_vector(0 to 31) := (others => '0');
    variable r2845 : std_logic_vector(0 to 31) := (others => '0');
    variable b2778 : boolean := false;
    variable r2777 : std_logic_vector(0 to 31) := (others => '0');
    variable r2776 : std_logic_vector(0 to 31) := (others => '0');
    variable b2709 : boolean := false;
    variable r2708 : std_logic_vector(0 to 31) := (others => '0');
    variable r2707 : std_logic_vector(0 to 31) := (others => '0');
    variable b2640 : boolean := false;
    variable r2639 : std_logic_vector(0 to 31) := (others => '0');
    variable r2638 : std_logic_vector(0 to 31) := (others => '0');
    variable b2571 : boolean := false;
    variable r2570 : std_logic_vector(0 to 31) := (others => '0');
    variable r2569 : std_logic_vector(0 to 31) := (others => '0');
    variable b2502 : boolean := false;
    variable r2501 : std_logic_vector(0 to 31) := (others => '0');
    variable r2500 : std_logic_vector(0 to 31) := (others => '0');
    variable b2433 : boolean := false;
    variable r2432 : std_logic_vector(0 to 31) := (others => '0');
    variable r2431 : std_logic_vector(0 to 31) := (others => '0');
    variable b2364 : boolean := false;
    variable r2363 : std_logic_vector(0 to 31) := (others => '0');
    variable r2362 : std_logic_vector(0 to 31) := (others => '0');
    variable b2295 : boolean := false;
    variable r2294 : std_logic_vector(0 to 31) := (others => '0');
    variable r2293 : std_logic_vector(0 to 31) := (others => '0');
    variable b2226 : boolean := false;
    variable r2225 : std_logic_vector(0 to 31) := (others => '0');
    variable r2224 : std_logic_vector(0 to 31) := (others => '0');
    variable b2157 : boolean := false;
    variable r2156 : std_logic_vector(0 to 31) := (others => '0');
    variable r2155 : std_logic_vector(0 to 31) := (others => '0');
    variable b2088 : boolean := false;
    variable r2087 : std_logic_vector(0 to 31) := (others => '0');
    variable r2086 : std_logic_vector(0 to 31) := (others => '0');
    variable b2019 : boolean := false;
    variable r2018 : std_logic_vector(0 to 31) := (others => '0');
    variable r2017 : std_logic_vector(0 to 31) := (others => '0');
    variable b1950 : boolean := false;
    variable r1949 : std_logic_vector(0 to 31) := (others => '0');
    variable r1948 : std_logic_vector(0 to 31) := (others => '0');
    variable b1881 : boolean := false;
    variable r1880 : std_logic_vector(0 to 31) := (others => '0');
    variable r1879 : std_logic_vector(0 to 31) := (others => '0');
    variable b1812 : boolean := false;
    variable r1811 : std_logic_vector(0 to 31) := (others => '0');
    variable r1810 : std_logic_vector(0 to 31) := (others => '0');
    variable b1743 : boolean := false;
    variable r1742 : std_logic_vector(0 to 31) := (others => '0');
    variable r1741 : std_logic_vector(0 to 31) := (others => '0');
    variable b1674 : boolean := false;
    variable r1673 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    b1674 := ("000000" = r1672(0 to 5));
    if b1674 then
      r1741 := rewire_MetaprogrammingRW.w428a2f98_1675;
      r1673 := r1741;
     else 
      null;
      b1743 := ("000001" = r1672(0 to 5));
      if b1743 then
        r1810 := rewire_MetaprogrammingRW.w71374491_1744;
        r1742 := r1810;
       else 
        null;
        b1812 := ("000010" = r1672(0 to 5));
        if b1812 then
          r1879 := rewire_MetaprogrammingRW.wb5c0fbcf_1813;
          r1811 := r1879;
         else 
          null;
          b1881 := ("000011" = r1672(0 to 5));
          if b1881 then
            r1948 := rewire_MetaprogrammingRW.we9b5dba5_1882;
            r1880 := r1948;
           else 
            null;
            b1950 := ("000100" = r1672(0 to 5));
            if b1950 then
              r2017 := rewire_MetaprogrammingRW.w3956c25b_1951;
              r1949 := r2017;
             else 
              null;
              b2019 := ("000101" = r1672(0 to 5));
              if b2019 then
                r2086 := rewire_MetaprogrammingRW.w59f111f1_2020;
                r2018 := r2086;
               else 
                null;
                b2088 := ("000110" = r1672(0 to 5));
                if b2088 then
                  r2155 := rewire_MetaprogrammingRW.w923f82a4_2089;
                  r2087 := r2155;
                 else 
                  null;
                  b2157 := ("000111" = r1672(0 to 5));
                  if b2157 then
                    r2224 := rewire_MetaprogrammingRW.wab1c5ed5_2158;
                    r2156 := r2224;
                   else 
                    null;
                    b2226 := ("001000" = r1672(0 to 5));
                    if b2226 then
                      r2293 := rewire_MetaprogrammingRW.wd807aa98_2227;
                      r2225 := r2293;
                     else 
                      null;
                      b2295 := ("001001" = r1672(0 to 5));
                      if b2295 then
                        r2362 := rewire_MetaprogrammingRW.w12835b01_2296;
                        r2294 := r2362;
                       else 
                        null;
                        b2364 := ("001010" = r1672(0 to 5));
                        if b2364 then
                          r2431 := rewire_MetaprogrammingRW.w243185be_2365;
                          r2363 := r2431;
                         else 
                          null;
                          b2433 := ("001011" = r1672(0 to 5));
                          if b2433 then
                            r2500 := rewire_MetaprogrammingRW.w550c7dc3_2434;
                            r2432 := r2500;
                           else 
                            null;
                            b2502 := ("001100" = r1672(0 to 5));
                            if b2502 then
                              r2569 := rewire_MetaprogrammingRW.w72be5d74_2503;
                              r2501 := r2569;
                             else 
                              null;
                              b2571 := ("001101" = r1672(0 to 5));
                              if b2571 then
                                r2638 := rewire_MetaprogrammingRW.w80deb1fe_2572;
                                r2570 := r2638;
                               else 
                                null;
                                b2640 := ("001110" = r1672(0 to 5));
                                if b2640 then
                                  r2707 := rewire_MetaprogrammingRW.w9bdc06a7_2641;
                                  r2639 := r2707;
                                 else 
                                  null;
                                  b2709 := ("001111" = r1672(0 to 5));
                                  if b2709 then
                                    r2776 := rewire_MetaprogrammingRW.wc19bf174_2710;
                                    r2708 := r2776;
                                   else 
                                    null;
                                    b2778 := ("010000" = r1672(0 to 5));
                                    if b2778 then
                                      r2845 := rewire_MetaprogrammingRW.we49b69c1_2779;
                                      r2777 := r2845;
                                     else 
                                      null;
                                      b2847 := ("010001" = r1672(0 to 5));
                                      if b2847 then
                                        r2914 := rewire_MetaprogrammingRW.wefbe4786_2848;
                                        r2846 := r2914;
                                       else 
                                        null;
                                        b2916 := ("010010" = r1672(0 to 5));
                                        if b2916 then
                                          r2983 := rewire_MetaprogrammingRW.w0fc19dc6_2917;
                                          r2915 := r2983;
                                         else 
                                          null;
                                          b2985 := ("010011" = r1672(0 to 5));
                                          if b2985 then
                                            r3052 := rewire_MetaprogrammingRW.w240ca1cc_2986;
                                            r2984 := r3052;
                                           else 
                                            null;
                                            b3054 := ("010100" = r1672(0 to 5));
                                            if b3054 then
                                              r3121 := rewire_MetaprogrammingRW.w2de92c6f_3055;
                                              r3053 := r3121;
                                             else 
                                              null;
                                              b3123 := ("010101" = r1672(0 to 5));
                                              if b3123 then
                                                r3190 := rewire_MetaprogrammingRW.w4a7484aa_3124;
                                                r3122 := r3190;
                                               else 
                                                null;
                                                b3192 := ("010110" = r1672(0 to 5));
                                                if b3192 then
                                                  r3259 := rewire_MetaprogrammingRW.w5cb0a9dc_3193;
                                                  r3191 := r3259;
                                                 else 
                                                  null;
                                                  b3261 := ("010111" = r1672(0 to 5));
                                                  if b3261 then
                                                    r3328 := rewire_MetaprogrammingRW.w76f988da_3262;
                                                    r3260 := r3328;
                                                   else 
                                                    null;
                                                    b3330 := ("011000" = r1672(0 to 5));
                                                    if b3330 then
                                                      r3397 := rewire_MetaprogrammingRW.w983e5152_3331;
                                                      r3329 := r3397;
                                                     else 
                                                      null;
                                                      b3399 := ("011001" = r1672(0 to 5));
                                                      if b3399 then
                                                        r3466 := rewire_MetaprogrammingRW.wa831c66d_3400;
                                                        r3398 := r3466;
                                                       else 
                                                        null;
                                                        b3468 := ("011010" = r1672(0 to 5));
                                                        if b3468 then
                                                          r3535 := rewire_MetaprogrammingRW.wb00327c8_3469;
                                                          r3467 := r3535;
                                                         else 
                                                          null;
                                                          b3537 := ("011011" = r1672(0 to 5));
                                                          if b3537 then
                                                            r3604 := rewire_MetaprogrammingRW.wbf597fc7_3538;
                                                            r3536 := r3604;
                                                           else 
                                                            null;
                                                            b3606 := ("011100" = r1672(0 to 5));
                                                            if b3606 then
                                                              r3673 := rewire_MetaprogrammingRW.wc6e00bf3_3607;
                                                              r3605 := r3673;
                                                             else 
                                                              null;
                                                              b3675 := ("011101" = r1672(0 to 5));
                                                              if b3675 then
                                                                r3742 := rewire_MetaprogrammingRW.wd5a79147_3676;
                                                                r3674 := r3742;
                                                               else 
                                                                null;
                                                                b3744 := ("011110" = r1672(0 to 5));
                                                                if b3744 then
                                                                  r3811 := rewire_MetaprogrammingRW.w06ca6351_3745;
                                                                  r3743 := r3811;
                                                                 else 
                                                                  null;
                                                                  b3813 := ("011111" = r1672(0 to 5));
                                                                  if b3813 then
                                                                    r3880 := rewire_MetaprogrammingRW.w14292967_3814;
                                                                    r3812 := r3880;
                                                                   else 
                                                                    null;
                                                                    b3882 := ("100000" = r1672(0 to 5));
                                                                    if b3882 then
                                                                      r3949 := rewire_MetaprogrammingRW.w27b70a85_3883;
                                                                      r3881 := r3949;
                                                                     else 
                                                                      null;
                                                                      b3951 := ("100001" = r1672(0 to 5));
                                                                      if b3951 then
                                                                        r4018 := rewire_MetaprogrammingRW.w2e1b2138_3952;
                                                                        r3950 := r4018;
                                                                       else 
                                                                        null;
                                                                        b4020 := ("100010" = r1672(0 to 5));
                                                                        if b4020 then
                                                                          r4087 := rewire_MetaprogrammingRW.w4d2c6dfc_4021;
                                                                          r4019 := r4087;
                                                                         else 
                                                                          null;
                                                                          b4089 := ("100011" = r1672(0 to 5));
                                                                          if b4089 then
                                                                            r4156 := rewire_MetaprogrammingRW.w53380d13_4090;
                                                                            r4088 := r4156;
                                                                           else 
                                                                            null;
                                                                            b4158 := ("100100" = r1672(0 to 5));
                                                                            if b4158 then
                                                                              r4225 := rewire_MetaprogrammingRW.w650a7354_4159;
                                                                              r4157 := r4225;
                                                                             else 
                                                                              null;
                                                                              b4227 := ("100101" = r1672(0 to 5));
                                                                              if b4227 then
                                                                                r4294 := rewire_MetaprogrammingRW.w766a0abb_4228;
                                                                                r4226 := r4294;
                                                                               else 
                                                                                null;
                                                                                b4296 := ("100110" = r1672(0 to 5));
                                                                                if b4296 then
                                                                                  r4363 := rewire_MetaprogrammingRW.w81c2c92e_4297;
                                                                                  r4295 := r4363;
                                                                                 else 
                                                                                  null;
                                                                                  b4365 := ("100111" = r1672(0 to 5));
                                                                                  if b4365 then
                                                                                    r4432 := rewire_MetaprogrammingRW.w92722c85_4366;
                                                                                    r4364 := r4432;
                                                                                   else 
                                                                                    null;
                                                                                    b4434 := ("101000" = r1672(0 to 5));
                                                                                    if b4434 then
                                                                                      r4501 := rewire_MetaprogrammingRW.wa2bfe8a1_4435;
                                                                                      r4433 := r4501;
                                                                                     else 
                                                                                      null;
                                                                                      b4503 := ("101001" = r1672(0 to 5));
                                                                                      if b4503 then
                                                                                        r4570 := rewire_MetaprogrammingRW.wa81a664b_4504;
                                                                                        r4502 := r4570;
                                                                                       else 
                                                                                        null;
                                                                                        b4572 := ("101010" = r1672(0 to 5));
                                                                                        if b4572 then
                                                                                          r4639 := rewire_MetaprogrammingRW.wc24b8b70_4573;
                                                                                          r4571 := r4639;
                                                                                         else 
                                                                                          null;
                                                                                          b4641 := ("101011" = r1672(0 to 5));
                                                                                          if b4641 then
                                                                                            r4708 := rewire_MetaprogrammingRW.wc76c51a3_4642;
                                                                                            r4640 := r4708;
                                                                                           else 
                                                                                            null;
                                                                                            b4710 := ("101100" = r1672(0 to 5));
                                                                                            if b4710 then
                                                                                              r4777 := rewire_MetaprogrammingRW.wd192e819_4711;
                                                                                              r4709 := r4777;
                                                                                             else 
                                                                                              null;
                                                                                              b4779 := ("101101" = r1672(0 to 5));
                                                                                              if b4779 then
                                                                                                r4846 := rewire_MetaprogrammingRW.wd6990624_4780;
                                                                                                r4778 := r4846;
                                                                                               else 
                                                                                                null;
                                                                                                b4848 := ("101110" = r1672(0 to 5));
                                                                                                if b4848 then
                                                                                                  r4915 := rewire_MetaprogrammingRW.wf40e3585_4849;
                                                                                                  r4847 := r4915;
                                                                                                 else 
                                                                                                  null;
                                                                                                  b4917 := ("101111" = r1672(0 to 5));
                                                                                                  if b4917 then
                                                                                                    r4984 := rewire_MetaprogrammingRW.w106aa070_4918;
                                                                                                    r4916 := r4984;
                                                                                                   else 
                                                                                                    null;
                                                                                                    b4986 := ("110000" = r1672(0 to 5));
                                                                                                    if b4986 then
                                                                                                      r5053 := rewire_MetaprogrammingRW.w19a4c116_4987;
                                                                                                      r4985 := r5053;
                                                                                                     else 
                                                                                                      null;
                                                                                                      b5055 := ("110001" = r1672(0 to 5));
                                                                                                      if b5055 then
                                                                                                        r5122 := rewire_MetaprogrammingRW.w1e376c08_5056;
                                                                                                        r5054 := r5122;
                                                                                                       else 
                                                                                                        null;
                                                                                                        b5124 := ("110010" = r1672(0 to 5));
                                                                                                        if b5124 then
                                                                                                          r5191 := rewire_MetaprogrammingRW.w2748774c_5125;
                                                                                                          r5123 := r5191;
                                                                                                         else 
                                                                                                          null;
                                                                                                          b5193 := ("110011" = r1672(0 to 5));
                                                                                                          if b5193 then
                                                                                                            r5260 := rewire_MetaprogrammingRW.w34b0bcb5_5194;
                                                                                                            r5192 := r5260;
                                                                                                           else 
                                                                                                            null;
                                                                                                            b5262 := ("110100" = r1672(0 to 5));
                                                                                                            if b5262 then
                                                                                                              r5329 := rewire_MetaprogrammingRW.w391c0cb3_5263;
                                                                                                              r5261 := r5329;
                                                                                                             else 
                                                                                                              null;
                                                                                                              b5331 := ("110101" = r1672(0 to 5));
                                                                                                              if b5331 then
                                                                                                                r5398 := rewire_MetaprogrammingRW.w4ed8aa4a_5332;
                                                                                                                r5330 := r5398;
                                                                                                               else 
                                                                                                                null;
                                                                                                                b5400 := ("110110" = r1672(0 to 5));
                                                                                                                if b5400 then
                                                                                                                  r5467 := rewire_MetaprogrammingRW.w5b9cca4f_5401;
                                                                                                                  r5399 := r5467;
                                                                                                                 else 
                                                                                                                  null;
                                                                                                                  b5469 := ("110111" = r1672(0 to 5));
                                                                                                                  if b5469 then
                                                                                                                    r5536 := rewire_MetaprogrammingRW.w682e6ff3_5470;
                                                                                                                    r5468 := r5536;
                                                                                                                   else 
                                                                                                                    null;
                                                                                                                    b5538 := ("111000" = r1672(0 to 5));
                                                                                                                    if b5538 then
                                                                                                                      r5605 := rewire_MetaprogrammingRW.w748f82ee_5539;
                                                                                                                      r5537 := r5605;
                                                                                                                     else 
                                                                                                                      null;
                                                                                                                      b5607 := ("111001" = r1672(0 to 5));
                                                                                                                      if b5607 then
                                                                                                                        r5674 := rewire_MetaprogrammingRW.w78a5636f_5608;
                                                                                                                        r5606 := r5674;
                                                                                                                       else 
                                                                                                                        null;
                                                                                                                        b5676 := ("111010" = r1672(0 to 5));
                                                                                                                        if b5676 then
                                                                                                                          r5743 := rewire_MetaprogrammingRW.w84c87814_5677;
                                                                                                                          r5675 := r5743;
                                                                                                                         else 
                                                                                                                          null;
                                                                                                                          b5745 := ("111011" = r1672(0 to 5));
                                                                                                                          if b5745 then
                                                                                                                            r5812 := rewire_MetaprogrammingRW.w8cc70208_5746;
                                                                                                                            r5744 := r5812;
                                                                                                                           else 
                                                                                                                            null;
                                                                                                                            b5814 := ("111100" = r1672(0 to 5));
                                                                                                                            if b5814 then
                                                                                                                              r5881 := rewire_MetaprogrammingRW.w90befffa_5815;
                                                                                                                              r5813 := r5881;
                                                                                                                             else 
                                                                                                                              null;
                                                                                                                              b5883 := ("111101" = r1672(0 to 5));
                                                                                                                              if b5883 then
                                                                                                                                r5950 := rewire_MetaprogrammingRW.wa4506ceb_5884;
                                                                                                                                r5882 := r5950;
                                                                                                                               else 
                                                                                                                                null;
                                                                                                                                b5952 := ("111110" = r1672(0 to 5));
                                                                                                                                if b5952 then
                                                                                                                                  r6019 := rewire_MetaprogrammingRW.wbef9a3f7_5953;
                                                                                                                                  r5951 := r6019;
                                                                                                                                 else 
                                                                                                                                  null;
                                                                                                                                  b6021 := ("111111" = r1672(0 to 5));
                                                                                                                                  r6088 := rewire_MetaprogrammingRW.wc67178f2_6022;
                                                                                                                                  r6020 := r6088;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;end if;
    return r1673;
  end rewire_Main.seed_1671;
  function rewire_MetaprogrammingRW.wc67178f2_6022 return std_logic_vector
  is
    variable r6087 : std_logic_vector(0 to 0) := (others => '0');
    variable r6086 : std_logic_vector(0 to 0) := (others => '0');
    variable r6085 : std_logic_vector(0 to 0) := (others => '0');
    variable r6084 : std_logic_vector(0 to 0) := (others => '0');
    variable r6083 : std_logic_vector(0 to 0) := (others => '0');
    variable r6082 : std_logic_vector(0 to 0) := (others => '0');
    variable r6081 : std_logic_vector(0 to 0) := (others => '0');
    variable r6080 : std_logic_vector(0 to 0) := (others => '0');
    variable r6079 : std_logic_vector(0 to 0) := (others => '0');
    variable r6078 : std_logic_vector(0 to 0) := (others => '0');
    variable r6077 : std_logic_vector(0 to 0) := (others => '0');
    variable r6076 : std_logic_vector(0 to 0) := (others => '0');
    variable r6075 : std_logic_vector(0 to 0) := (others => '0');
    variable r6074 : std_logic_vector(0 to 0) := (others => '0');
    variable r6073 : std_logic_vector(0 to 0) := (others => '0');
    variable r6072 : std_logic_vector(0 to 0) := (others => '0');
    variable r6071 : std_logic_vector(0 to 0) := (others => '0');
    variable r6070 : std_logic_vector(0 to 0) := (others => '0');
    variable r6069 : std_logic_vector(0 to 0) := (others => '0');
    variable r6068 : std_logic_vector(0 to 0) := (others => '0');
    variable r6067 : std_logic_vector(0 to 0) := (others => '0');
    variable r6066 : std_logic_vector(0 to 0) := (others => '0');
    variable r6065 : std_logic_vector(0 to 0) := (others => '0');
    variable r6064 : std_logic_vector(0 to 0) := (others => '0');
    variable r6063 : std_logic_vector(0 to 0) := (others => '0');
    variable r6062 : std_logic_vector(0 to 0) := (others => '0');
    variable r6061 : std_logic_vector(0 to 0) := (others => '0');
    variable r6060 : std_logic_vector(0 to 0) := (others => '0');
    variable r6059 : std_logic_vector(0 to 0) := (others => '0');
    variable r6058 : std_logic_vector(0 to 0) := (others => '0');
    variable r6057 : std_logic_vector(0 to 0) := (others => '0');
    variable r6056 : std_logic_vector(0 to 0) := (others => '0');
    variable r6055 : std_logic_vector(0 to 0) := (others => '0');
    variable r6054 : std_logic_vector(0 to 0) := (others => '0');
    variable r6053 : std_logic_vector(0 to 0) := (others => '0');
    variable r6052 : std_logic_vector(0 to 0) := (others => '0');
    variable r6051 : std_logic_vector(0 to 0) := (others => '0');
    variable r6050 : std_logic_vector(0 to 0) := (others => '0');
    variable r6049 : std_logic_vector(0 to 0) := (others => '0');
    variable r6048 : std_logic_vector(0 to 0) := (others => '0');
    variable r6047 : std_logic_vector(0 to 0) := (others => '0');
    variable r6046 : std_logic_vector(0 to 0) := (others => '0');
    variable r6045 : std_logic_vector(0 to 0) := (others => '0');
    variable r6044 : std_logic_vector(0 to 0) := (others => '0');
    variable r6043 : std_logic_vector(0 to 0) := (others => '0');
    variable r6042 : std_logic_vector(0 to 0) := (others => '0');
    variable r6041 : std_logic_vector(0 to 0) := (others => '0');
    variable r6040 : std_logic_vector(0 to 0) := (others => '0');
    variable r6039 : std_logic_vector(0 to 0) := (others => '0');
    variable r6038 : std_logic_vector(0 to 0) := (others => '0');
    variable r6037 : std_logic_vector(0 to 0) := (others => '0');
    variable r6036 : std_logic_vector(0 to 0) := (others => '0');
    variable r6035 : std_logic_vector(0 to 0) := (others => '0');
    variable r6034 : std_logic_vector(0 to 0) := (others => '0');
    variable r6033 : std_logic_vector(0 to 0) := (others => '0');
    variable r6032 : std_logic_vector(0 to 0) := (others => '0');
    variable r6031 : std_logic_vector(0 to 0) := (others => '0');
    variable r6030 : std_logic_vector(0 to 0) := (others => '0');
    variable r6029 : std_logic_vector(0 to 0) := (others => '0');
    variable r6028 : std_logic_vector(0 to 0) := (others => '0');
    variable r6027 : std_logic_vector(0 to 0) := (others => '0');
    variable r6026 : std_logic_vector(0 to 0) := (others => '0');
    variable r6025 : std_logic_vector(0 to 0) := (others => '0');
    variable r6024 : std_logic_vector(0 to 0) := (others => '0');
    variable r6023 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r6024 := "1";
    null;
    r6025 := (r6024);
    r6026 := "1";
    null;
    r6027 := (r6026);
    r6028 := "0";
    null;
    r6029 := (r6028);
    r6030 := "0";
    null;
    r6031 := (r6030);
    r6032 := "0";
    null;
    r6033 := (r6032);
    r6034 := "1";
    null;
    r6035 := (r6034);
    r6036 := "1";
    null;
    r6037 := (r6036);
    r6038 := "0";
    null;
    r6039 := (r6038);
    r6040 := "0";
    null;
    r6041 := (r6040);
    r6042 := "1";
    null;
    r6043 := (r6042);
    r6044 := "1";
    null;
    r6045 := (r6044);
    r6046 := "1";
    null;
    r6047 := (r6046);
    r6048 := "0";
    null;
    r6049 := (r6048);
    r6050 := "0";
    null;
    r6051 := (r6050);
    r6052 := "0";
    null;
    r6053 := (r6052);
    r6054 := "1";
    null;
    r6055 := (r6054);
    r6056 := "0";
    null;
    r6057 := (r6056);
    r6058 := "1";
    null;
    r6059 := (r6058);
    r6060 := "1";
    null;
    r6061 := (r6060);
    r6062 := "1";
    null;
    r6063 := (r6062);
    r6064 := "1";
    null;
    r6065 := (r6064);
    r6066 := "0";
    null;
    r6067 := (r6066);
    r6068 := "0";
    null;
    r6069 := (r6068);
    r6070 := "0";
    null;
    r6071 := (r6070);
    r6072 := "1";
    null;
    r6073 := (r6072);
    r6074 := "1";
    null;
    r6075 := (r6074);
    r6076 := "1";
    null;
    r6077 := (r6076);
    r6078 := "1";
    null;
    r6079 := (r6078);
    r6080 := "0";
    null;
    r6081 := (r6080);
    r6082 := "0";
    null;
    r6083 := (r6082);
    r6084 := "1";
    null;
    r6085 := (r6084);
    r6086 := "0";
    null;
    r6087 := (r6086);
    r6023 := (r6025 & r6027 & r6029 & r6031 & r6033 & r6035 & r6037 & r6039 & r6041 & r6043 & r6045 & r6047 & r6049 & r6051 & r6053 & r6055 & r6057 & r6059 & r6061 & r6063 & r6065 & r6067 & r6069 & r6071 & r6073 & r6075 & r6077 & r6079 & r6081 & r6083 & r6085 & r6087);
    return r6023;
  end rewire_MetaprogrammingRW.wc67178f2_6022;
  function rewire_MetaprogrammingRW.wbef9a3f7_5953 return std_logic_vector
  is
    variable r6018 : std_logic_vector(0 to 0) := (others => '0');
    variable r6017 : std_logic_vector(0 to 0) := (others => '0');
    variable r6016 : std_logic_vector(0 to 0) := (others => '0');
    variable r6015 : std_logic_vector(0 to 0) := (others => '0');
    variable r6014 : std_logic_vector(0 to 0) := (others => '0');
    variable r6013 : std_logic_vector(0 to 0) := (others => '0');
    variable r6012 : std_logic_vector(0 to 0) := (others => '0');
    variable r6011 : std_logic_vector(0 to 0) := (others => '0');
    variable r6010 : std_logic_vector(0 to 0) := (others => '0');
    variable r6009 : std_logic_vector(0 to 0) := (others => '0');
    variable r6008 : std_logic_vector(0 to 0) := (others => '0');
    variable r6007 : std_logic_vector(0 to 0) := (others => '0');
    variable r6006 : std_logic_vector(0 to 0) := (others => '0');
    variable r6005 : std_logic_vector(0 to 0) := (others => '0');
    variable r6004 : std_logic_vector(0 to 0) := (others => '0');
    variable r6003 : std_logic_vector(0 to 0) := (others => '0');
    variable r6002 : std_logic_vector(0 to 0) := (others => '0');
    variable r6001 : std_logic_vector(0 to 0) := (others => '0');
    variable r6000 : std_logic_vector(0 to 0) := (others => '0');
    variable r5999 : std_logic_vector(0 to 0) := (others => '0');
    variable r5998 : std_logic_vector(0 to 0) := (others => '0');
    variable r5997 : std_logic_vector(0 to 0) := (others => '0');
    variable r5996 : std_logic_vector(0 to 0) := (others => '0');
    variable r5995 : std_logic_vector(0 to 0) := (others => '0');
    variable r5994 : std_logic_vector(0 to 0) := (others => '0');
    variable r5993 : std_logic_vector(0 to 0) := (others => '0');
    variable r5992 : std_logic_vector(0 to 0) := (others => '0');
    variable r5991 : std_logic_vector(0 to 0) := (others => '0');
    variable r5990 : std_logic_vector(0 to 0) := (others => '0');
    variable r5989 : std_logic_vector(0 to 0) := (others => '0');
    variable r5988 : std_logic_vector(0 to 0) := (others => '0');
    variable r5987 : std_logic_vector(0 to 0) := (others => '0');
    variable r5986 : std_logic_vector(0 to 0) := (others => '0');
    variable r5985 : std_logic_vector(0 to 0) := (others => '0');
    variable r5984 : std_logic_vector(0 to 0) := (others => '0');
    variable r5983 : std_logic_vector(0 to 0) := (others => '0');
    variable r5982 : std_logic_vector(0 to 0) := (others => '0');
    variable r5981 : std_logic_vector(0 to 0) := (others => '0');
    variable r5980 : std_logic_vector(0 to 0) := (others => '0');
    variable r5979 : std_logic_vector(0 to 0) := (others => '0');
    variable r5978 : std_logic_vector(0 to 0) := (others => '0');
    variable r5977 : std_logic_vector(0 to 0) := (others => '0');
    variable r5976 : std_logic_vector(0 to 0) := (others => '0');
    variable r5975 : std_logic_vector(0 to 0) := (others => '0');
    variable r5974 : std_logic_vector(0 to 0) := (others => '0');
    variable r5973 : std_logic_vector(0 to 0) := (others => '0');
    variable r5972 : std_logic_vector(0 to 0) := (others => '0');
    variable r5971 : std_logic_vector(0 to 0) := (others => '0');
    variable r5970 : std_logic_vector(0 to 0) := (others => '0');
    variable r5969 : std_logic_vector(0 to 0) := (others => '0');
    variable r5968 : std_logic_vector(0 to 0) := (others => '0');
    variable r5967 : std_logic_vector(0 to 0) := (others => '0');
    variable r5966 : std_logic_vector(0 to 0) := (others => '0');
    variable r5965 : std_logic_vector(0 to 0) := (others => '0');
    variable r5964 : std_logic_vector(0 to 0) := (others => '0');
    variable r5963 : std_logic_vector(0 to 0) := (others => '0');
    variable r5962 : std_logic_vector(0 to 0) := (others => '0');
    variable r5961 : std_logic_vector(0 to 0) := (others => '0');
    variable r5960 : std_logic_vector(0 to 0) := (others => '0');
    variable r5959 : std_logic_vector(0 to 0) := (others => '0');
    variable r5958 : std_logic_vector(0 to 0) := (others => '0');
    variable r5957 : std_logic_vector(0 to 0) := (others => '0');
    variable r5956 : std_logic_vector(0 to 0) := (others => '0');
    variable r5955 : std_logic_vector(0 to 0) := (others => '0');
    variable r5954 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r5955 := "1";
    null;
    r5956 := (r5955);
    r5957 := "0";
    null;
    r5958 := (r5957);
    r5959 := "1";
    null;
    r5960 := (r5959);
    r5961 := "1";
    null;
    r5962 := (r5961);
    r5963 := "1";
    null;
    r5964 := (r5963);
    r5965 := "1";
    null;
    r5966 := (r5965);
    r5967 := "1";
    null;
    r5968 := (r5967);
    r5969 := "0";
    null;
    r5970 := (r5969);
    r5971 := "1";
    null;
    r5972 := (r5971);
    r5973 := "1";
    null;
    r5974 := (r5973);
    r5975 := "1";
    null;
    r5976 := (r5975);
    r5977 := "1";
    null;
    r5978 := (r5977);
    r5979 := "1";
    null;
    r5980 := (r5979);
    r5981 := "0";
    null;
    r5982 := (r5981);
    r5983 := "0";
    null;
    r5984 := (r5983);
    r5985 := "1";
    null;
    r5986 := (r5985);
    r5987 := "1";
    null;
    r5988 := (r5987);
    r5989 := "0";
    null;
    r5990 := (r5989);
    r5991 := "1";
    null;
    r5992 := (r5991);
    r5993 := "0";
    null;
    r5994 := (r5993);
    r5995 := "0";
    null;
    r5996 := (r5995);
    r5997 := "0";
    null;
    r5998 := (r5997);
    r5999 := "1";
    null;
    r6000 := (r5999);
    r6001 := "1";
    null;
    r6002 := (r6001);
    r6003 := "1";
    null;
    r6004 := (r6003);
    r6005 := "1";
    null;
    r6006 := (r6005);
    r6007 := "1";
    null;
    r6008 := (r6007);
    r6009 := "1";
    null;
    r6010 := (r6009);
    r6011 := "0";
    null;
    r6012 := (r6011);
    r6013 := "1";
    null;
    r6014 := (r6013);
    r6015 := "1";
    null;
    r6016 := (r6015);
    r6017 := "1";
    null;
    r6018 := (r6017);
    r5954 := (r5956 & r5958 & r5960 & r5962 & r5964 & r5966 & r5968 & r5970 & r5972 & r5974 & r5976 & r5978 & r5980 & r5982 & r5984 & r5986 & r5988 & r5990 & r5992 & r5994 & r5996 & r5998 & r6000 & r6002 & r6004 & r6006 & r6008 & r6010 & r6012 & r6014 & r6016 & r6018);
    return r5954;
  end rewire_MetaprogrammingRW.wbef9a3f7_5953;
  function rewire_MetaprogrammingRW.wa4506ceb_5884 return std_logic_vector
  is
    variable r5949 : std_logic_vector(0 to 0) := (others => '0');
    variable r5948 : std_logic_vector(0 to 0) := (others => '0');
    variable r5947 : std_logic_vector(0 to 0) := (others => '0');
    variable r5946 : std_logic_vector(0 to 0) := (others => '0');
    variable r5945 : std_logic_vector(0 to 0) := (others => '0');
    variable r5944 : std_logic_vector(0 to 0) := (others => '0');
    variable r5943 : std_logic_vector(0 to 0) := (others => '0');
    variable r5942 : std_logic_vector(0 to 0) := (others => '0');
    variable r5941 : std_logic_vector(0 to 0) := (others => '0');
    variable r5940 : std_logic_vector(0 to 0) := (others => '0');
    variable r5939 : std_logic_vector(0 to 0) := (others => '0');
    variable r5938 : std_logic_vector(0 to 0) := (others => '0');
    variable r5937 : std_logic_vector(0 to 0) := (others => '0');
    variable r5936 : std_logic_vector(0 to 0) := (others => '0');
    variable r5935 : std_logic_vector(0 to 0) := (others => '0');
    variable r5934 : std_logic_vector(0 to 0) := (others => '0');
    variable r5933 : std_logic_vector(0 to 0) := (others => '0');
    variable r5932 : std_logic_vector(0 to 0) := (others => '0');
    variable r5931 : std_logic_vector(0 to 0) := (others => '0');
    variable r5930 : std_logic_vector(0 to 0) := (others => '0');
    variable r5929 : std_logic_vector(0 to 0) := (others => '0');
    variable r5928 : std_logic_vector(0 to 0) := (others => '0');
    variable r5927 : std_logic_vector(0 to 0) := (others => '0');
    variable r5926 : std_logic_vector(0 to 0) := (others => '0');
    variable r5925 : std_logic_vector(0 to 0) := (others => '0');
    variable r5924 : std_logic_vector(0 to 0) := (others => '0');
    variable r5923 : std_logic_vector(0 to 0) := (others => '0');
    variable r5922 : std_logic_vector(0 to 0) := (others => '0');
    variable r5921 : std_logic_vector(0 to 0) := (others => '0');
    variable r5920 : std_logic_vector(0 to 0) := (others => '0');
    variable r5919 : std_logic_vector(0 to 0) := (others => '0');
    variable r5918 : std_logic_vector(0 to 0) := (others => '0');
    variable r5917 : std_logic_vector(0 to 0) := (others => '0');
    variable r5916 : std_logic_vector(0 to 0) := (others => '0');
    variable r5915 : std_logic_vector(0 to 0) := (others => '0');
    variable r5914 : std_logic_vector(0 to 0) := (others => '0');
    variable r5913 : std_logic_vector(0 to 0) := (others => '0');
    variable r5912 : std_logic_vector(0 to 0) := (others => '0');
    variable r5911 : std_logic_vector(0 to 0) := (others => '0');
    variable r5910 : std_logic_vector(0 to 0) := (others => '0');
    variable r5909 : std_logic_vector(0 to 0) := (others => '0');
    variable r5908 : std_logic_vector(0 to 0) := (others => '0');
    variable r5907 : std_logic_vector(0 to 0) := (others => '0');
    variable r5906 : std_logic_vector(0 to 0) := (others => '0');
    variable r5905 : std_logic_vector(0 to 0) := (others => '0');
    variable r5904 : std_logic_vector(0 to 0) := (others => '0');
    variable r5903 : std_logic_vector(0 to 0) := (others => '0');
    variable r5902 : std_logic_vector(0 to 0) := (others => '0');
    variable r5901 : std_logic_vector(0 to 0) := (others => '0');
    variable r5900 : std_logic_vector(0 to 0) := (others => '0');
    variable r5899 : std_logic_vector(0 to 0) := (others => '0');
    variable r5898 : std_logic_vector(0 to 0) := (others => '0');
    variable r5897 : std_logic_vector(0 to 0) := (others => '0');
    variable r5896 : std_logic_vector(0 to 0) := (others => '0');
    variable r5895 : std_logic_vector(0 to 0) := (others => '0');
    variable r5894 : std_logic_vector(0 to 0) := (others => '0');
    variable r5893 : std_logic_vector(0 to 0) := (others => '0');
    variable r5892 : std_logic_vector(0 to 0) := (others => '0');
    variable r5891 : std_logic_vector(0 to 0) := (others => '0');
    variable r5890 : std_logic_vector(0 to 0) := (others => '0');
    variable r5889 : std_logic_vector(0 to 0) := (others => '0');
    variable r5888 : std_logic_vector(0 to 0) := (others => '0');
    variable r5887 : std_logic_vector(0 to 0) := (others => '0');
    variable r5886 : std_logic_vector(0 to 0) := (others => '0');
    variable r5885 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r5886 := "1";
    null;
    r5887 := (r5886);
    r5888 := "0";
    null;
    r5889 := (r5888);
    r5890 := "1";
    null;
    r5891 := (r5890);
    r5892 := "0";
    null;
    r5893 := (r5892);
    r5894 := "0";
    null;
    r5895 := (r5894);
    r5896 := "1";
    null;
    r5897 := (r5896);
    r5898 := "0";
    null;
    r5899 := (r5898);
    r5900 := "0";
    null;
    r5901 := (r5900);
    r5902 := "0";
    null;
    r5903 := (r5902);
    r5904 := "1";
    null;
    r5905 := (r5904);
    r5906 := "0";
    null;
    r5907 := (r5906);
    r5908 := "1";
    null;
    r5909 := (r5908);
    r5910 := "0";
    null;
    r5911 := (r5910);
    r5912 := "0";
    null;
    r5913 := (r5912);
    r5914 := "0";
    null;
    r5915 := (r5914);
    r5916 := "0";
    null;
    r5917 := (r5916);
    r5918 := "0";
    null;
    r5919 := (r5918);
    r5920 := "1";
    null;
    r5921 := (r5920);
    r5922 := "1";
    null;
    r5923 := (r5922);
    r5924 := "0";
    null;
    r5925 := (r5924);
    r5926 := "1";
    null;
    r5927 := (r5926);
    r5928 := "1";
    null;
    r5929 := (r5928);
    r5930 := "0";
    null;
    r5931 := (r5930);
    r5932 := "0";
    null;
    r5933 := (r5932);
    r5934 := "1";
    null;
    r5935 := (r5934);
    r5936 := "1";
    null;
    r5937 := (r5936);
    r5938 := "1";
    null;
    r5939 := (r5938);
    r5940 := "0";
    null;
    r5941 := (r5940);
    r5942 := "1";
    null;
    r5943 := (r5942);
    r5944 := "0";
    null;
    r5945 := (r5944);
    r5946 := "1";
    null;
    r5947 := (r5946);
    r5948 := "1";
    null;
    r5949 := (r5948);
    r5885 := (r5887 & r5889 & r5891 & r5893 & r5895 & r5897 & r5899 & r5901 & r5903 & r5905 & r5907 & r5909 & r5911 & r5913 & r5915 & r5917 & r5919 & r5921 & r5923 & r5925 & r5927 & r5929 & r5931 & r5933 & r5935 & r5937 & r5939 & r5941 & r5943 & r5945 & r5947 & r5949);
    return r5885;
  end rewire_MetaprogrammingRW.wa4506ceb_5884;
  function rewire_MetaprogrammingRW.w90befffa_5815 return std_logic_vector
  is
    variable r5880 : std_logic_vector(0 to 0) := (others => '0');
    variable r5879 : std_logic_vector(0 to 0) := (others => '0');
    variable r5878 : std_logic_vector(0 to 0) := (others => '0');
    variable r5877 : std_logic_vector(0 to 0) := (others => '0');
    variable r5876 : std_logic_vector(0 to 0) := (others => '0');
    variable r5875 : std_logic_vector(0 to 0) := (others => '0');
    variable r5874 : std_logic_vector(0 to 0) := (others => '0');
    variable r5873 : std_logic_vector(0 to 0) := (others => '0');
    variable r5872 : std_logic_vector(0 to 0) := (others => '0');
    variable r5871 : std_logic_vector(0 to 0) := (others => '0');
    variable r5870 : std_logic_vector(0 to 0) := (others => '0');
    variable r5869 : std_logic_vector(0 to 0) := (others => '0');
    variable r5868 : std_logic_vector(0 to 0) := (others => '0');
    variable r5867 : std_logic_vector(0 to 0) := (others => '0');
    variable r5866 : std_logic_vector(0 to 0) := (others => '0');
    variable r5865 : std_logic_vector(0 to 0) := (others => '0');
    variable r5864 : std_logic_vector(0 to 0) := (others => '0');
    variable r5863 : std_logic_vector(0 to 0) := (others => '0');
    variable r5862 : std_logic_vector(0 to 0) := (others => '0');
    variable r5861 : std_logic_vector(0 to 0) := (others => '0');
    variable r5860 : std_logic_vector(0 to 0) := (others => '0');
    variable r5859 : std_logic_vector(0 to 0) := (others => '0');
    variable r5858 : std_logic_vector(0 to 0) := (others => '0');
    variable r5857 : std_logic_vector(0 to 0) := (others => '0');
    variable r5856 : std_logic_vector(0 to 0) := (others => '0');
    variable r5855 : std_logic_vector(0 to 0) := (others => '0');
    variable r5854 : std_logic_vector(0 to 0) := (others => '0');
    variable r5853 : std_logic_vector(0 to 0) := (others => '0');
    variable r5852 : std_logic_vector(0 to 0) := (others => '0');
    variable r5851 : std_logic_vector(0 to 0) := (others => '0');
    variable r5850 : std_logic_vector(0 to 0) := (others => '0');
    variable r5849 : std_logic_vector(0 to 0) := (others => '0');
    variable r5848 : std_logic_vector(0 to 0) := (others => '0');
    variable r5847 : std_logic_vector(0 to 0) := (others => '0');
    variable r5846 : std_logic_vector(0 to 0) := (others => '0');
    variable r5845 : std_logic_vector(0 to 0) := (others => '0');
    variable r5844 : std_logic_vector(0 to 0) := (others => '0');
    variable r5843 : std_logic_vector(0 to 0) := (others => '0');
    variable r5842 : std_logic_vector(0 to 0) := (others => '0');
    variable r5841 : std_logic_vector(0 to 0) := (others => '0');
    variable r5840 : std_logic_vector(0 to 0) := (others => '0');
    variable r5839 : std_logic_vector(0 to 0) := (others => '0');
    variable r5838 : std_logic_vector(0 to 0) := (others => '0');
    variable r5837 : std_logic_vector(0 to 0) := (others => '0');
    variable r5836 : std_logic_vector(0 to 0) := (others => '0');
    variable r5835 : std_logic_vector(0 to 0) := (others => '0');
    variable r5834 : std_logic_vector(0 to 0) := (others => '0');
    variable r5833 : std_logic_vector(0 to 0) := (others => '0');
    variable r5832 : std_logic_vector(0 to 0) := (others => '0');
    variable r5831 : std_logic_vector(0 to 0) := (others => '0');
    variable r5830 : std_logic_vector(0 to 0) := (others => '0');
    variable r5829 : std_logic_vector(0 to 0) := (others => '0');
    variable r5828 : std_logic_vector(0 to 0) := (others => '0');
    variable r5827 : std_logic_vector(0 to 0) := (others => '0');
    variable r5826 : std_logic_vector(0 to 0) := (others => '0');
    variable r5825 : std_logic_vector(0 to 0) := (others => '0');
    variable r5824 : std_logic_vector(0 to 0) := (others => '0');
    variable r5823 : std_logic_vector(0 to 0) := (others => '0');
    variable r5822 : std_logic_vector(0 to 0) := (others => '0');
    variable r5821 : std_logic_vector(0 to 0) := (others => '0');
    variable r5820 : std_logic_vector(0 to 0) := (others => '0');
    variable r5819 : std_logic_vector(0 to 0) := (others => '0');
    variable r5818 : std_logic_vector(0 to 0) := (others => '0');
    variable r5817 : std_logic_vector(0 to 0) := (others => '0');
    variable r5816 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r5817 := "1";
    null;
    r5818 := (r5817);
    r5819 := "0";
    null;
    r5820 := (r5819);
    r5821 := "0";
    null;
    r5822 := (r5821);
    r5823 := "1";
    null;
    r5824 := (r5823);
    r5825 := "0";
    null;
    r5826 := (r5825);
    r5827 := "0";
    null;
    r5828 := (r5827);
    r5829 := "0";
    null;
    r5830 := (r5829);
    r5831 := "0";
    null;
    r5832 := (r5831);
    r5833 := "1";
    null;
    r5834 := (r5833);
    r5835 := "0";
    null;
    r5836 := (r5835);
    r5837 := "1";
    null;
    r5838 := (r5837);
    r5839 := "1";
    null;
    r5840 := (r5839);
    r5841 := "1";
    null;
    r5842 := (r5841);
    r5843 := "1";
    null;
    r5844 := (r5843);
    r5845 := "1";
    null;
    r5846 := (r5845);
    r5847 := "0";
    null;
    r5848 := (r5847);
    r5849 := "1";
    null;
    r5850 := (r5849);
    r5851 := "1";
    null;
    r5852 := (r5851);
    r5853 := "1";
    null;
    r5854 := (r5853);
    r5855 := "1";
    null;
    r5856 := (r5855);
    r5857 := "1";
    null;
    r5858 := (r5857);
    r5859 := "1";
    null;
    r5860 := (r5859);
    r5861 := "1";
    null;
    r5862 := (r5861);
    r5863 := "1";
    null;
    r5864 := (r5863);
    r5865 := "1";
    null;
    r5866 := (r5865);
    r5867 := "1";
    null;
    r5868 := (r5867);
    r5869 := "1";
    null;
    r5870 := (r5869);
    r5871 := "1";
    null;
    r5872 := (r5871);
    r5873 := "1";
    null;
    r5874 := (r5873);
    r5875 := "0";
    null;
    r5876 := (r5875);
    r5877 := "1";
    null;
    r5878 := (r5877);
    r5879 := "0";
    null;
    r5880 := (r5879);
    r5816 := (r5818 & r5820 & r5822 & r5824 & r5826 & r5828 & r5830 & r5832 & r5834 & r5836 & r5838 & r5840 & r5842 & r5844 & r5846 & r5848 & r5850 & r5852 & r5854 & r5856 & r5858 & r5860 & r5862 & r5864 & r5866 & r5868 & r5870 & r5872 & r5874 & r5876 & r5878 & r5880);
    return r5816;
  end rewire_MetaprogrammingRW.w90befffa_5815;
  function rewire_MetaprogrammingRW.w8cc70208_5746 return std_logic_vector
  is
    variable r5811 : std_logic_vector(0 to 0) := (others => '0');
    variable r5810 : std_logic_vector(0 to 0) := (others => '0');
    variable r5809 : std_logic_vector(0 to 0) := (others => '0');
    variable r5808 : std_logic_vector(0 to 0) := (others => '0');
    variable r5807 : std_logic_vector(0 to 0) := (others => '0');
    variable r5806 : std_logic_vector(0 to 0) := (others => '0');
    variable r5805 : std_logic_vector(0 to 0) := (others => '0');
    variable r5804 : std_logic_vector(0 to 0) := (others => '0');
    variable r5803 : std_logic_vector(0 to 0) := (others => '0');
    variable r5802 : std_logic_vector(0 to 0) := (others => '0');
    variable r5801 : std_logic_vector(0 to 0) := (others => '0');
    variable r5800 : std_logic_vector(0 to 0) := (others => '0');
    variable r5799 : std_logic_vector(0 to 0) := (others => '0');
    variable r5798 : std_logic_vector(0 to 0) := (others => '0');
    variable r5797 : std_logic_vector(0 to 0) := (others => '0');
    variable r5796 : std_logic_vector(0 to 0) := (others => '0');
    variable r5795 : std_logic_vector(0 to 0) := (others => '0');
    variable r5794 : std_logic_vector(0 to 0) := (others => '0');
    variable r5793 : std_logic_vector(0 to 0) := (others => '0');
    variable r5792 : std_logic_vector(0 to 0) := (others => '0');
    variable r5791 : std_logic_vector(0 to 0) := (others => '0');
    variable r5790 : std_logic_vector(0 to 0) := (others => '0');
    variable r5789 : std_logic_vector(0 to 0) := (others => '0');
    variable r5788 : std_logic_vector(0 to 0) := (others => '0');
    variable r5787 : std_logic_vector(0 to 0) := (others => '0');
    variable r5786 : std_logic_vector(0 to 0) := (others => '0');
    variable r5785 : std_logic_vector(0 to 0) := (others => '0');
    variable r5784 : std_logic_vector(0 to 0) := (others => '0');
    variable r5783 : std_logic_vector(0 to 0) := (others => '0');
    variable r5782 : std_logic_vector(0 to 0) := (others => '0');
    variable r5781 : std_logic_vector(0 to 0) := (others => '0');
    variable r5780 : std_logic_vector(0 to 0) := (others => '0');
    variable r5779 : std_logic_vector(0 to 0) := (others => '0');
    variable r5778 : std_logic_vector(0 to 0) := (others => '0');
    variable r5777 : std_logic_vector(0 to 0) := (others => '0');
    variable r5776 : std_logic_vector(0 to 0) := (others => '0');
    variable r5775 : std_logic_vector(0 to 0) := (others => '0');
    variable r5774 : std_logic_vector(0 to 0) := (others => '0');
    variable r5773 : std_logic_vector(0 to 0) := (others => '0');
    variable r5772 : std_logic_vector(0 to 0) := (others => '0');
    variable r5771 : std_logic_vector(0 to 0) := (others => '0');
    variable r5770 : std_logic_vector(0 to 0) := (others => '0');
    variable r5769 : std_logic_vector(0 to 0) := (others => '0');
    variable r5768 : std_logic_vector(0 to 0) := (others => '0');
    variable r5767 : std_logic_vector(0 to 0) := (others => '0');
    variable r5766 : std_logic_vector(0 to 0) := (others => '0');
    variable r5765 : std_logic_vector(0 to 0) := (others => '0');
    variable r5764 : std_logic_vector(0 to 0) := (others => '0');
    variable r5763 : std_logic_vector(0 to 0) := (others => '0');
    variable r5762 : std_logic_vector(0 to 0) := (others => '0');
    variable r5761 : std_logic_vector(0 to 0) := (others => '0');
    variable r5760 : std_logic_vector(0 to 0) := (others => '0');
    variable r5759 : std_logic_vector(0 to 0) := (others => '0');
    variable r5758 : std_logic_vector(0 to 0) := (others => '0');
    variable r5757 : std_logic_vector(0 to 0) := (others => '0');
    variable r5756 : std_logic_vector(0 to 0) := (others => '0');
    variable r5755 : std_logic_vector(0 to 0) := (others => '0');
    variable r5754 : std_logic_vector(0 to 0) := (others => '0');
    variable r5753 : std_logic_vector(0 to 0) := (others => '0');
    variable r5752 : std_logic_vector(0 to 0) := (others => '0');
    variable r5751 : std_logic_vector(0 to 0) := (others => '0');
    variable r5750 : std_logic_vector(0 to 0) := (others => '0');
    variable r5749 : std_logic_vector(0 to 0) := (others => '0');
    variable r5748 : std_logic_vector(0 to 0) := (others => '0');
    variable r5747 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r5748 := "1";
    null;
    r5749 := (r5748);
    r5750 := "0";
    null;
    r5751 := (r5750);
    r5752 := "0";
    null;
    r5753 := (r5752);
    r5754 := "0";
    null;
    r5755 := (r5754);
    r5756 := "1";
    null;
    r5757 := (r5756);
    r5758 := "1";
    null;
    r5759 := (r5758);
    r5760 := "0";
    null;
    r5761 := (r5760);
    r5762 := "0";
    null;
    r5763 := (r5762);
    r5764 := "1";
    null;
    r5765 := (r5764);
    r5766 := "1";
    null;
    r5767 := (r5766);
    r5768 := "0";
    null;
    r5769 := (r5768);
    r5770 := "0";
    null;
    r5771 := (r5770);
    r5772 := "0";
    null;
    r5773 := (r5772);
    r5774 := "1";
    null;
    r5775 := (r5774);
    r5776 := "1";
    null;
    r5777 := (r5776);
    r5778 := "1";
    null;
    r5779 := (r5778);
    r5780 := "0";
    null;
    r5781 := (r5780);
    r5782 := "0";
    null;
    r5783 := (r5782);
    r5784 := "0";
    null;
    r5785 := (r5784);
    r5786 := "0";
    null;
    r5787 := (r5786);
    r5788 := "0";
    null;
    r5789 := (r5788);
    r5790 := "0";
    null;
    r5791 := (r5790);
    r5792 := "1";
    null;
    r5793 := (r5792);
    r5794 := "0";
    null;
    r5795 := (r5794);
    r5796 := "0";
    null;
    r5797 := (r5796);
    r5798 := "0";
    null;
    r5799 := (r5798);
    r5800 := "0";
    null;
    r5801 := (r5800);
    r5802 := "0";
    null;
    r5803 := (r5802);
    r5804 := "1";
    null;
    r5805 := (r5804);
    r5806 := "0";
    null;
    r5807 := (r5806);
    r5808 := "0";
    null;
    r5809 := (r5808);
    r5810 := "0";
    null;
    r5811 := (r5810);
    r5747 := (r5749 & r5751 & r5753 & r5755 & r5757 & r5759 & r5761 & r5763 & r5765 & r5767 & r5769 & r5771 & r5773 & r5775 & r5777 & r5779 & r5781 & r5783 & r5785 & r5787 & r5789 & r5791 & r5793 & r5795 & r5797 & r5799 & r5801 & r5803 & r5805 & r5807 & r5809 & r5811);
    return r5747;
  end rewire_MetaprogrammingRW.w8cc70208_5746;
  function rewire_MetaprogrammingRW.w84c87814_5677 return std_logic_vector
  is
    variable r5742 : std_logic_vector(0 to 0) := (others => '0');
    variable r5741 : std_logic_vector(0 to 0) := (others => '0');
    variable r5740 : std_logic_vector(0 to 0) := (others => '0');
    variable r5739 : std_logic_vector(0 to 0) := (others => '0');
    variable r5738 : std_logic_vector(0 to 0) := (others => '0');
    variable r5737 : std_logic_vector(0 to 0) := (others => '0');
    variable r5736 : std_logic_vector(0 to 0) := (others => '0');
    variable r5735 : std_logic_vector(0 to 0) := (others => '0');
    variable r5734 : std_logic_vector(0 to 0) := (others => '0');
    variable r5733 : std_logic_vector(0 to 0) := (others => '0');
    variable r5732 : std_logic_vector(0 to 0) := (others => '0');
    variable r5731 : std_logic_vector(0 to 0) := (others => '0');
    variable r5730 : std_logic_vector(0 to 0) := (others => '0');
    variable r5729 : std_logic_vector(0 to 0) := (others => '0');
    variable r5728 : std_logic_vector(0 to 0) := (others => '0');
    variable r5727 : std_logic_vector(0 to 0) := (others => '0');
    variable r5726 : std_logic_vector(0 to 0) := (others => '0');
    variable r5725 : std_logic_vector(0 to 0) := (others => '0');
    variable r5724 : std_logic_vector(0 to 0) := (others => '0');
    variable r5723 : std_logic_vector(0 to 0) := (others => '0');
    variable r5722 : std_logic_vector(0 to 0) := (others => '0');
    variable r5721 : std_logic_vector(0 to 0) := (others => '0');
    variable r5720 : std_logic_vector(0 to 0) := (others => '0');
    variable r5719 : std_logic_vector(0 to 0) := (others => '0');
    variable r5718 : std_logic_vector(0 to 0) := (others => '0');
    variable r5717 : std_logic_vector(0 to 0) := (others => '0');
    variable r5716 : std_logic_vector(0 to 0) := (others => '0');
    variable r5715 : std_logic_vector(0 to 0) := (others => '0');
    variable r5714 : std_logic_vector(0 to 0) := (others => '0');
    variable r5713 : std_logic_vector(0 to 0) := (others => '0');
    variable r5712 : std_logic_vector(0 to 0) := (others => '0');
    variable r5711 : std_logic_vector(0 to 0) := (others => '0');
    variable r5710 : std_logic_vector(0 to 0) := (others => '0');
    variable r5709 : std_logic_vector(0 to 0) := (others => '0');
    variable r5708 : std_logic_vector(0 to 0) := (others => '0');
    variable r5707 : std_logic_vector(0 to 0) := (others => '0');
    variable r5706 : std_logic_vector(0 to 0) := (others => '0');
    variable r5705 : std_logic_vector(0 to 0) := (others => '0');
    variable r5704 : std_logic_vector(0 to 0) := (others => '0');
    variable r5703 : std_logic_vector(0 to 0) := (others => '0');
    variable r5702 : std_logic_vector(0 to 0) := (others => '0');
    variable r5701 : std_logic_vector(0 to 0) := (others => '0');
    variable r5700 : std_logic_vector(0 to 0) := (others => '0');
    variable r5699 : std_logic_vector(0 to 0) := (others => '0');
    variable r5698 : std_logic_vector(0 to 0) := (others => '0');
    variable r5697 : std_logic_vector(0 to 0) := (others => '0');
    variable r5696 : std_logic_vector(0 to 0) := (others => '0');
    variable r5695 : std_logic_vector(0 to 0) := (others => '0');
    variable r5694 : std_logic_vector(0 to 0) := (others => '0');
    variable r5693 : std_logic_vector(0 to 0) := (others => '0');
    variable r5692 : std_logic_vector(0 to 0) := (others => '0');
    variable r5691 : std_logic_vector(0 to 0) := (others => '0');
    variable r5690 : std_logic_vector(0 to 0) := (others => '0');
    variable r5689 : std_logic_vector(0 to 0) := (others => '0');
    variable r5688 : std_logic_vector(0 to 0) := (others => '0');
    variable r5687 : std_logic_vector(0 to 0) := (others => '0');
    variable r5686 : std_logic_vector(0 to 0) := (others => '0');
    variable r5685 : std_logic_vector(0 to 0) := (others => '0');
    variable r5684 : std_logic_vector(0 to 0) := (others => '0');
    variable r5683 : std_logic_vector(0 to 0) := (others => '0');
    variable r5682 : std_logic_vector(0 to 0) := (others => '0');
    variable r5681 : std_logic_vector(0 to 0) := (others => '0');
    variable r5680 : std_logic_vector(0 to 0) := (others => '0');
    variable r5679 : std_logic_vector(0 to 0) := (others => '0');
    variable r5678 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r5679 := "1";
    null;
    r5680 := (r5679);
    r5681 := "0";
    null;
    r5682 := (r5681);
    r5683 := "0";
    null;
    r5684 := (r5683);
    r5685 := "0";
    null;
    r5686 := (r5685);
    r5687 := "0";
    null;
    r5688 := (r5687);
    r5689 := "1";
    null;
    r5690 := (r5689);
    r5691 := "0";
    null;
    r5692 := (r5691);
    r5693 := "0";
    null;
    r5694 := (r5693);
    r5695 := "1";
    null;
    r5696 := (r5695);
    r5697 := "1";
    null;
    r5698 := (r5697);
    r5699 := "0";
    null;
    r5700 := (r5699);
    r5701 := "0";
    null;
    r5702 := (r5701);
    r5703 := "1";
    null;
    r5704 := (r5703);
    r5705 := "0";
    null;
    r5706 := (r5705);
    r5707 := "0";
    null;
    r5708 := (r5707);
    r5709 := "0";
    null;
    r5710 := (r5709);
    r5711 := "0";
    null;
    r5712 := (r5711);
    r5713 := "1";
    null;
    r5714 := (r5713);
    r5715 := "1";
    null;
    r5716 := (r5715);
    r5717 := "1";
    null;
    r5718 := (r5717);
    r5719 := "1";
    null;
    r5720 := (r5719);
    r5721 := "0";
    null;
    r5722 := (r5721);
    r5723 := "0";
    null;
    r5724 := (r5723);
    r5725 := "0";
    null;
    r5726 := (r5725);
    r5727 := "0";
    null;
    r5728 := (r5727);
    r5729 := "0";
    null;
    r5730 := (r5729);
    r5731 := "0";
    null;
    r5732 := (r5731);
    r5733 := "1";
    null;
    r5734 := (r5733);
    r5735 := "0";
    null;
    r5736 := (r5735);
    r5737 := "1";
    null;
    r5738 := (r5737);
    r5739 := "0";
    null;
    r5740 := (r5739);
    r5741 := "0";
    null;
    r5742 := (r5741);
    r5678 := (r5680 & r5682 & r5684 & r5686 & r5688 & r5690 & r5692 & r5694 & r5696 & r5698 & r5700 & r5702 & r5704 & r5706 & r5708 & r5710 & r5712 & r5714 & r5716 & r5718 & r5720 & r5722 & r5724 & r5726 & r5728 & r5730 & r5732 & r5734 & r5736 & r5738 & r5740 & r5742);
    return r5678;
  end rewire_MetaprogrammingRW.w84c87814_5677;
  function rewire_MetaprogrammingRW.w78a5636f_5608 return std_logic_vector
  is
    variable r5673 : std_logic_vector(0 to 0) := (others => '0');
    variable r5672 : std_logic_vector(0 to 0) := (others => '0');
    variable r5671 : std_logic_vector(0 to 0) := (others => '0');
    variable r5670 : std_logic_vector(0 to 0) := (others => '0');
    variable r5669 : std_logic_vector(0 to 0) := (others => '0');
    variable r5668 : std_logic_vector(0 to 0) := (others => '0');
    variable r5667 : std_logic_vector(0 to 0) := (others => '0');
    variable r5666 : std_logic_vector(0 to 0) := (others => '0');
    variable r5665 : std_logic_vector(0 to 0) := (others => '0');
    variable r5664 : std_logic_vector(0 to 0) := (others => '0');
    variable r5663 : std_logic_vector(0 to 0) := (others => '0');
    variable r5662 : std_logic_vector(0 to 0) := (others => '0');
    variable r5661 : std_logic_vector(0 to 0) := (others => '0');
    variable r5660 : std_logic_vector(0 to 0) := (others => '0');
    variable r5659 : std_logic_vector(0 to 0) := (others => '0');
    variable r5658 : std_logic_vector(0 to 0) := (others => '0');
    variable r5657 : std_logic_vector(0 to 0) := (others => '0');
    variable r5656 : std_logic_vector(0 to 0) := (others => '0');
    variable r5655 : std_logic_vector(0 to 0) := (others => '0');
    variable r5654 : std_logic_vector(0 to 0) := (others => '0');
    variable r5653 : std_logic_vector(0 to 0) := (others => '0');
    variable r5652 : std_logic_vector(0 to 0) := (others => '0');
    variable r5651 : std_logic_vector(0 to 0) := (others => '0');
    variable r5650 : std_logic_vector(0 to 0) := (others => '0');
    variable r5649 : std_logic_vector(0 to 0) := (others => '0');
    variable r5648 : std_logic_vector(0 to 0) := (others => '0');
    variable r5647 : std_logic_vector(0 to 0) := (others => '0');
    variable r5646 : std_logic_vector(0 to 0) := (others => '0');
    variable r5645 : std_logic_vector(0 to 0) := (others => '0');
    variable r5644 : std_logic_vector(0 to 0) := (others => '0');
    variable r5643 : std_logic_vector(0 to 0) := (others => '0');
    variable r5642 : std_logic_vector(0 to 0) := (others => '0');
    variable r5641 : std_logic_vector(0 to 0) := (others => '0');
    variable r5640 : std_logic_vector(0 to 0) := (others => '0');
    variable r5639 : std_logic_vector(0 to 0) := (others => '0');
    variable r5638 : std_logic_vector(0 to 0) := (others => '0');
    variable r5637 : std_logic_vector(0 to 0) := (others => '0');
    variable r5636 : std_logic_vector(0 to 0) := (others => '0');
    variable r5635 : std_logic_vector(0 to 0) := (others => '0');
    variable r5634 : std_logic_vector(0 to 0) := (others => '0');
    variable r5633 : std_logic_vector(0 to 0) := (others => '0');
    variable r5632 : std_logic_vector(0 to 0) := (others => '0');
    variable r5631 : std_logic_vector(0 to 0) := (others => '0');
    variable r5630 : std_logic_vector(0 to 0) := (others => '0');
    variable r5629 : std_logic_vector(0 to 0) := (others => '0');
    variable r5628 : std_logic_vector(0 to 0) := (others => '0');
    variable r5627 : std_logic_vector(0 to 0) := (others => '0');
    variable r5626 : std_logic_vector(0 to 0) := (others => '0');
    variable r5625 : std_logic_vector(0 to 0) := (others => '0');
    variable r5624 : std_logic_vector(0 to 0) := (others => '0');
    variable r5623 : std_logic_vector(0 to 0) := (others => '0');
    variable r5622 : std_logic_vector(0 to 0) := (others => '0');
    variable r5621 : std_logic_vector(0 to 0) := (others => '0');
    variable r5620 : std_logic_vector(0 to 0) := (others => '0');
    variable r5619 : std_logic_vector(0 to 0) := (others => '0');
    variable r5618 : std_logic_vector(0 to 0) := (others => '0');
    variable r5617 : std_logic_vector(0 to 0) := (others => '0');
    variable r5616 : std_logic_vector(0 to 0) := (others => '0');
    variable r5615 : std_logic_vector(0 to 0) := (others => '0');
    variable r5614 : std_logic_vector(0 to 0) := (others => '0');
    variable r5613 : std_logic_vector(0 to 0) := (others => '0');
    variable r5612 : std_logic_vector(0 to 0) := (others => '0');
    variable r5611 : std_logic_vector(0 to 0) := (others => '0');
    variable r5610 : std_logic_vector(0 to 0) := (others => '0');
    variable r5609 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r5610 := "0";
    null;
    r5611 := (r5610);
    r5612 := "1";
    null;
    r5613 := (r5612);
    r5614 := "1";
    null;
    r5615 := (r5614);
    r5616 := "1";
    null;
    r5617 := (r5616);
    r5618 := "1";
    null;
    r5619 := (r5618);
    r5620 := "0";
    null;
    r5621 := (r5620);
    r5622 := "0";
    null;
    r5623 := (r5622);
    r5624 := "0";
    null;
    r5625 := (r5624);
    r5626 := "1";
    null;
    r5627 := (r5626);
    r5628 := "0";
    null;
    r5629 := (r5628);
    r5630 := "1";
    null;
    r5631 := (r5630);
    r5632 := "0";
    null;
    r5633 := (r5632);
    r5634 := "0";
    null;
    r5635 := (r5634);
    r5636 := "1";
    null;
    r5637 := (r5636);
    r5638 := "0";
    null;
    r5639 := (r5638);
    r5640 := "1";
    null;
    r5641 := (r5640);
    r5642 := "0";
    null;
    r5643 := (r5642);
    r5644 := "1";
    null;
    r5645 := (r5644);
    r5646 := "1";
    null;
    r5647 := (r5646);
    r5648 := "0";
    null;
    r5649 := (r5648);
    r5650 := "0";
    null;
    r5651 := (r5650);
    r5652 := "0";
    null;
    r5653 := (r5652);
    r5654 := "1";
    null;
    r5655 := (r5654);
    r5656 := "1";
    null;
    r5657 := (r5656);
    r5658 := "0";
    null;
    r5659 := (r5658);
    r5660 := "1";
    null;
    r5661 := (r5660);
    r5662 := "1";
    null;
    r5663 := (r5662);
    r5664 := "0";
    null;
    r5665 := (r5664);
    r5666 := "1";
    null;
    r5667 := (r5666);
    r5668 := "1";
    null;
    r5669 := (r5668);
    r5670 := "1";
    null;
    r5671 := (r5670);
    r5672 := "1";
    null;
    r5673 := (r5672);
    r5609 := (r5611 & r5613 & r5615 & r5617 & r5619 & r5621 & r5623 & r5625 & r5627 & r5629 & r5631 & r5633 & r5635 & r5637 & r5639 & r5641 & r5643 & r5645 & r5647 & r5649 & r5651 & r5653 & r5655 & r5657 & r5659 & r5661 & r5663 & r5665 & r5667 & r5669 & r5671 & r5673);
    return r5609;
  end rewire_MetaprogrammingRW.w78a5636f_5608;
  function rewire_MetaprogrammingRW.w748f82ee_5539 return std_logic_vector
  is
    variable r5604 : std_logic_vector(0 to 0) := (others => '0');
    variable r5603 : std_logic_vector(0 to 0) := (others => '0');
    variable r5602 : std_logic_vector(0 to 0) := (others => '0');
    variable r5601 : std_logic_vector(0 to 0) := (others => '0');
    variable r5600 : std_logic_vector(0 to 0) := (others => '0');
    variable r5599 : std_logic_vector(0 to 0) := (others => '0');
    variable r5598 : std_logic_vector(0 to 0) := (others => '0');
    variable r5597 : std_logic_vector(0 to 0) := (others => '0');
    variable r5596 : std_logic_vector(0 to 0) := (others => '0');
    variable r5595 : std_logic_vector(0 to 0) := (others => '0');
    variable r5594 : std_logic_vector(0 to 0) := (others => '0');
    variable r5593 : std_logic_vector(0 to 0) := (others => '0');
    variable r5592 : std_logic_vector(0 to 0) := (others => '0');
    variable r5591 : std_logic_vector(0 to 0) := (others => '0');
    variable r5590 : std_logic_vector(0 to 0) := (others => '0');
    variable r5589 : std_logic_vector(0 to 0) := (others => '0');
    variable r5588 : std_logic_vector(0 to 0) := (others => '0');
    variable r5587 : std_logic_vector(0 to 0) := (others => '0');
    variable r5586 : std_logic_vector(0 to 0) := (others => '0');
    variable r5585 : std_logic_vector(0 to 0) := (others => '0');
    variable r5584 : std_logic_vector(0 to 0) := (others => '0');
    variable r5583 : std_logic_vector(0 to 0) := (others => '0');
    variable r5582 : std_logic_vector(0 to 0) := (others => '0');
    variable r5581 : std_logic_vector(0 to 0) := (others => '0');
    variable r5580 : std_logic_vector(0 to 0) := (others => '0');
    variable r5579 : std_logic_vector(0 to 0) := (others => '0');
    variable r5578 : std_logic_vector(0 to 0) := (others => '0');
    variable r5577 : std_logic_vector(0 to 0) := (others => '0');
    variable r5576 : std_logic_vector(0 to 0) := (others => '0');
    variable r5575 : std_logic_vector(0 to 0) := (others => '0');
    variable r5574 : std_logic_vector(0 to 0) := (others => '0');
    variable r5573 : std_logic_vector(0 to 0) := (others => '0');
    variable r5572 : std_logic_vector(0 to 0) := (others => '0');
    variable r5571 : std_logic_vector(0 to 0) := (others => '0');
    variable r5570 : std_logic_vector(0 to 0) := (others => '0');
    variable r5569 : std_logic_vector(0 to 0) := (others => '0');
    variable r5568 : std_logic_vector(0 to 0) := (others => '0');
    variable r5567 : std_logic_vector(0 to 0) := (others => '0');
    variable r5566 : std_logic_vector(0 to 0) := (others => '0');
    variable r5565 : std_logic_vector(0 to 0) := (others => '0');
    variable r5564 : std_logic_vector(0 to 0) := (others => '0');
    variable r5563 : std_logic_vector(0 to 0) := (others => '0');
    variable r5562 : std_logic_vector(0 to 0) := (others => '0');
    variable r5561 : std_logic_vector(0 to 0) := (others => '0');
    variable r5560 : std_logic_vector(0 to 0) := (others => '0');
    variable r5559 : std_logic_vector(0 to 0) := (others => '0');
    variable r5558 : std_logic_vector(0 to 0) := (others => '0');
    variable r5557 : std_logic_vector(0 to 0) := (others => '0');
    variable r5556 : std_logic_vector(0 to 0) := (others => '0');
    variable r5555 : std_logic_vector(0 to 0) := (others => '0');
    variable r5554 : std_logic_vector(0 to 0) := (others => '0');
    variable r5553 : std_logic_vector(0 to 0) := (others => '0');
    variable r5552 : std_logic_vector(0 to 0) := (others => '0');
    variable r5551 : std_logic_vector(0 to 0) := (others => '0');
    variable r5550 : std_logic_vector(0 to 0) := (others => '0');
    variable r5549 : std_logic_vector(0 to 0) := (others => '0');
    variable r5548 : std_logic_vector(0 to 0) := (others => '0');
    variable r5547 : std_logic_vector(0 to 0) := (others => '0');
    variable r5546 : std_logic_vector(0 to 0) := (others => '0');
    variable r5545 : std_logic_vector(0 to 0) := (others => '0');
    variable r5544 : std_logic_vector(0 to 0) := (others => '0');
    variable r5543 : std_logic_vector(0 to 0) := (others => '0');
    variable r5542 : std_logic_vector(0 to 0) := (others => '0');
    variable r5541 : std_logic_vector(0 to 0) := (others => '0');
    variable r5540 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r5541 := "0";
    null;
    r5542 := (r5541);
    r5543 := "1";
    null;
    r5544 := (r5543);
    r5545 := "1";
    null;
    r5546 := (r5545);
    r5547 := "1";
    null;
    r5548 := (r5547);
    r5549 := "0";
    null;
    r5550 := (r5549);
    r5551 := "1";
    null;
    r5552 := (r5551);
    r5553 := "0";
    null;
    r5554 := (r5553);
    r5555 := "0";
    null;
    r5556 := (r5555);
    r5557 := "1";
    null;
    r5558 := (r5557);
    r5559 := "0";
    null;
    r5560 := (r5559);
    r5561 := "0";
    null;
    r5562 := (r5561);
    r5563 := "0";
    null;
    r5564 := (r5563);
    r5565 := "1";
    null;
    r5566 := (r5565);
    r5567 := "1";
    null;
    r5568 := (r5567);
    r5569 := "1";
    null;
    r5570 := (r5569);
    r5571 := "1";
    null;
    r5572 := (r5571);
    r5573 := "1";
    null;
    r5574 := (r5573);
    r5575 := "0";
    null;
    r5576 := (r5575);
    r5577 := "0";
    null;
    r5578 := (r5577);
    r5579 := "0";
    null;
    r5580 := (r5579);
    r5581 := "0";
    null;
    r5582 := (r5581);
    r5583 := "0";
    null;
    r5584 := (r5583);
    r5585 := "1";
    null;
    r5586 := (r5585);
    r5587 := "0";
    null;
    r5588 := (r5587);
    r5589 := "1";
    null;
    r5590 := (r5589);
    r5591 := "1";
    null;
    r5592 := (r5591);
    r5593 := "1";
    null;
    r5594 := (r5593);
    r5595 := "0";
    null;
    r5596 := (r5595);
    r5597 := "1";
    null;
    r5598 := (r5597);
    r5599 := "1";
    null;
    r5600 := (r5599);
    r5601 := "1";
    null;
    r5602 := (r5601);
    r5603 := "0";
    null;
    r5604 := (r5603);
    r5540 := (r5542 & r5544 & r5546 & r5548 & r5550 & r5552 & r5554 & r5556 & r5558 & r5560 & r5562 & r5564 & r5566 & r5568 & r5570 & r5572 & r5574 & r5576 & r5578 & r5580 & r5582 & r5584 & r5586 & r5588 & r5590 & r5592 & r5594 & r5596 & r5598 & r5600 & r5602 & r5604);
    return r5540;
  end rewire_MetaprogrammingRW.w748f82ee_5539;
  function rewire_MetaprogrammingRW.w682e6ff3_5470 return std_logic_vector
  is
    variable r5535 : std_logic_vector(0 to 0) := (others => '0');
    variable r5534 : std_logic_vector(0 to 0) := (others => '0');
    variable r5533 : std_logic_vector(0 to 0) := (others => '0');
    variable r5532 : std_logic_vector(0 to 0) := (others => '0');
    variable r5531 : std_logic_vector(0 to 0) := (others => '0');
    variable r5530 : std_logic_vector(0 to 0) := (others => '0');
    variable r5529 : std_logic_vector(0 to 0) := (others => '0');
    variable r5528 : std_logic_vector(0 to 0) := (others => '0');
    variable r5527 : std_logic_vector(0 to 0) := (others => '0');
    variable r5526 : std_logic_vector(0 to 0) := (others => '0');
    variable r5525 : std_logic_vector(0 to 0) := (others => '0');
    variable r5524 : std_logic_vector(0 to 0) := (others => '0');
    variable r5523 : std_logic_vector(0 to 0) := (others => '0');
    variable r5522 : std_logic_vector(0 to 0) := (others => '0');
    variable r5521 : std_logic_vector(0 to 0) := (others => '0');
    variable r5520 : std_logic_vector(0 to 0) := (others => '0');
    variable r5519 : std_logic_vector(0 to 0) := (others => '0');
    variable r5518 : std_logic_vector(0 to 0) := (others => '0');
    variable r5517 : std_logic_vector(0 to 0) := (others => '0');
    variable r5516 : std_logic_vector(0 to 0) := (others => '0');
    variable r5515 : std_logic_vector(0 to 0) := (others => '0');
    variable r5514 : std_logic_vector(0 to 0) := (others => '0');
    variable r5513 : std_logic_vector(0 to 0) := (others => '0');
    variable r5512 : std_logic_vector(0 to 0) := (others => '0');
    variable r5511 : std_logic_vector(0 to 0) := (others => '0');
    variable r5510 : std_logic_vector(0 to 0) := (others => '0');
    variable r5509 : std_logic_vector(0 to 0) := (others => '0');
    variable r5508 : std_logic_vector(0 to 0) := (others => '0');
    variable r5507 : std_logic_vector(0 to 0) := (others => '0');
    variable r5506 : std_logic_vector(0 to 0) := (others => '0');
    variable r5505 : std_logic_vector(0 to 0) := (others => '0');
    variable r5504 : std_logic_vector(0 to 0) := (others => '0');
    variable r5503 : std_logic_vector(0 to 0) := (others => '0');
    variable r5502 : std_logic_vector(0 to 0) := (others => '0');
    variable r5501 : std_logic_vector(0 to 0) := (others => '0');
    variable r5500 : std_logic_vector(0 to 0) := (others => '0');
    variable r5499 : std_logic_vector(0 to 0) := (others => '0');
    variable r5498 : std_logic_vector(0 to 0) := (others => '0');
    variable r5497 : std_logic_vector(0 to 0) := (others => '0');
    variable r5496 : std_logic_vector(0 to 0) := (others => '0');
    variable r5495 : std_logic_vector(0 to 0) := (others => '0');
    variable r5494 : std_logic_vector(0 to 0) := (others => '0');
    variable r5493 : std_logic_vector(0 to 0) := (others => '0');
    variable r5492 : std_logic_vector(0 to 0) := (others => '0');
    variable r5491 : std_logic_vector(0 to 0) := (others => '0');
    variable r5490 : std_logic_vector(0 to 0) := (others => '0');
    variable r5489 : std_logic_vector(0 to 0) := (others => '0');
    variable r5488 : std_logic_vector(0 to 0) := (others => '0');
    variable r5487 : std_logic_vector(0 to 0) := (others => '0');
    variable r5486 : std_logic_vector(0 to 0) := (others => '0');
    variable r5485 : std_logic_vector(0 to 0) := (others => '0');
    variable r5484 : std_logic_vector(0 to 0) := (others => '0');
    variable r5483 : std_logic_vector(0 to 0) := (others => '0');
    variable r5482 : std_logic_vector(0 to 0) := (others => '0');
    variable r5481 : std_logic_vector(0 to 0) := (others => '0');
    variable r5480 : std_logic_vector(0 to 0) := (others => '0');
    variable r5479 : std_logic_vector(0 to 0) := (others => '0');
    variable r5478 : std_logic_vector(0 to 0) := (others => '0');
    variable r5477 : std_logic_vector(0 to 0) := (others => '0');
    variable r5476 : std_logic_vector(0 to 0) := (others => '0');
    variable r5475 : std_logic_vector(0 to 0) := (others => '0');
    variable r5474 : std_logic_vector(0 to 0) := (others => '0');
    variable r5473 : std_logic_vector(0 to 0) := (others => '0');
    variable r5472 : std_logic_vector(0 to 0) := (others => '0');
    variable r5471 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r5472 := "0";
    null;
    r5473 := (r5472);
    r5474 := "1";
    null;
    r5475 := (r5474);
    r5476 := "1";
    null;
    r5477 := (r5476);
    r5478 := "0";
    null;
    r5479 := (r5478);
    r5480 := "1";
    null;
    r5481 := (r5480);
    r5482 := "0";
    null;
    r5483 := (r5482);
    r5484 := "0";
    null;
    r5485 := (r5484);
    r5486 := "0";
    null;
    r5487 := (r5486);
    r5488 := "0";
    null;
    r5489 := (r5488);
    r5490 := "0";
    null;
    r5491 := (r5490);
    r5492 := "1";
    null;
    r5493 := (r5492);
    r5494 := "0";
    null;
    r5495 := (r5494);
    r5496 := "1";
    null;
    r5497 := (r5496);
    r5498 := "1";
    null;
    r5499 := (r5498);
    r5500 := "1";
    null;
    r5501 := (r5500);
    r5502 := "0";
    null;
    r5503 := (r5502);
    r5504 := "0";
    null;
    r5505 := (r5504);
    r5506 := "1";
    null;
    r5507 := (r5506);
    r5508 := "1";
    null;
    r5509 := (r5508);
    r5510 := "0";
    null;
    r5511 := (r5510);
    r5512 := "1";
    null;
    r5513 := (r5512);
    r5514 := "1";
    null;
    r5515 := (r5514);
    r5516 := "1";
    null;
    r5517 := (r5516);
    r5518 := "1";
    null;
    r5519 := (r5518);
    r5520 := "1";
    null;
    r5521 := (r5520);
    r5522 := "1";
    null;
    r5523 := (r5522);
    r5524 := "1";
    null;
    r5525 := (r5524);
    r5526 := "1";
    null;
    r5527 := (r5526);
    r5528 := "0";
    null;
    r5529 := (r5528);
    r5530 := "0";
    null;
    r5531 := (r5530);
    r5532 := "1";
    null;
    r5533 := (r5532);
    r5534 := "1";
    null;
    r5535 := (r5534);
    r5471 := (r5473 & r5475 & r5477 & r5479 & r5481 & r5483 & r5485 & r5487 & r5489 & r5491 & r5493 & r5495 & r5497 & r5499 & r5501 & r5503 & r5505 & r5507 & r5509 & r5511 & r5513 & r5515 & r5517 & r5519 & r5521 & r5523 & r5525 & r5527 & r5529 & r5531 & r5533 & r5535);
    return r5471;
  end rewire_MetaprogrammingRW.w682e6ff3_5470;
  function rewire_MetaprogrammingRW.w5b9cca4f_5401 return std_logic_vector
  is
    variable r5466 : std_logic_vector(0 to 0) := (others => '0');
    variable r5465 : std_logic_vector(0 to 0) := (others => '0');
    variable r5464 : std_logic_vector(0 to 0) := (others => '0');
    variable r5463 : std_logic_vector(0 to 0) := (others => '0');
    variable r5462 : std_logic_vector(0 to 0) := (others => '0');
    variable r5461 : std_logic_vector(0 to 0) := (others => '0');
    variable r5460 : std_logic_vector(0 to 0) := (others => '0');
    variable r5459 : std_logic_vector(0 to 0) := (others => '0');
    variable r5458 : std_logic_vector(0 to 0) := (others => '0');
    variable r5457 : std_logic_vector(0 to 0) := (others => '0');
    variable r5456 : std_logic_vector(0 to 0) := (others => '0');
    variable r5455 : std_logic_vector(0 to 0) := (others => '0');
    variable r5454 : std_logic_vector(0 to 0) := (others => '0');
    variable r5453 : std_logic_vector(0 to 0) := (others => '0');
    variable r5452 : std_logic_vector(0 to 0) := (others => '0');
    variable r5451 : std_logic_vector(0 to 0) := (others => '0');
    variable r5450 : std_logic_vector(0 to 0) := (others => '0');
    variable r5449 : std_logic_vector(0 to 0) := (others => '0');
    variable r5448 : std_logic_vector(0 to 0) := (others => '0');
    variable r5447 : std_logic_vector(0 to 0) := (others => '0');
    variable r5446 : std_logic_vector(0 to 0) := (others => '0');
    variable r5445 : std_logic_vector(0 to 0) := (others => '0');
    variable r5444 : std_logic_vector(0 to 0) := (others => '0');
    variable r5443 : std_logic_vector(0 to 0) := (others => '0');
    variable r5442 : std_logic_vector(0 to 0) := (others => '0');
    variable r5441 : std_logic_vector(0 to 0) := (others => '0');
    variable r5440 : std_logic_vector(0 to 0) := (others => '0');
    variable r5439 : std_logic_vector(0 to 0) := (others => '0');
    variable r5438 : std_logic_vector(0 to 0) := (others => '0');
    variable r5437 : std_logic_vector(0 to 0) := (others => '0');
    variable r5436 : std_logic_vector(0 to 0) := (others => '0');
    variable r5435 : std_logic_vector(0 to 0) := (others => '0');
    variable r5434 : std_logic_vector(0 to 0) := (others => '0');
    variable r5433 : std_logic_vector(0 to 0) := (others => '0');
    variable r5432 : std_logic_vector(0 to 0) := (others => '0');
    variable r5431 : std_logic_vector(0 to 0) := (others => '0');
    variable r5430 : std_logic_vector(0 to 0) := (others => '0');
    variable r5429 : std_logic_vector(0 to 0) := (others => '0');
    variable r5428 : std_logic_vector(0 to 0) := (others => '0');
    variable r5427 : std_logic_vector(0 to 0) := (others => '0');
    variable r5426 : std_logic_vector(0 to 0) := (others => '0');
    variable r5425 : std_logic_vector(0 to 0) := (others => '0');
    variable r5424 : std_logic_vector(0 to 0) := (others => '0');
    variable r5423 : std_logic_vector(0 to 0) := (others => '0');
    variable r5422 : std_logic_vector(0 to 0) := (others => '0');
    variable r5421 : std_logic_vector(0 to 0) := (others => '0');
    variable r5420 : std_logic_vector(0 to 0) := (others => '0');
    variable r5419 : std_logic_vector(0 to 0) := (others => '0');
    variable r5418 : std_logic_vector(0 to 0) := (others => '0');
    variable r5417 : std_logic_vector(0 to 0) := (others => '0');
    variable r5416 : std_logic_vector(0 to 0) := (others => '0');
    variable r5415 : std_logic_vector(0 to 0) := (others => '0');
    variable r5414 : std_logic_vector(0 to 0) := (others => '0');
    variable r5413 : std_logic_vector(0 to 0) := (others => '0');
    variable r5412 : std_logic_vector(0 to 0) := (others => '0');
    variable r5411 : std_logic_vector(0 to 0) := (others => '0');
    variable r5410 : std_logic_vector(0 to 0) := (others => '0');
    variable r5409 : std_logic_vector(0 to 0) := (others => '0');
    variable r5408 : std_logic_vector(0 to 0) := (others => '0');
    variable r5407 : std_logic_vector(0 to 0) := (others => '0');
    variable r5406 : std_logic_vector(0 to 0) := (others => '0');
    variable r5405 : std_logic_vector(0 to 0) := (others => '0');
    variable r5404 : std_logic_vector(0 to 0) := (others => '0');
    variable r5403 : std_logic_vector(0 to 0) := (others => '0');
    variable r5402 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r5403 := "0";
    null;
    r5404 := (r5403);
    r5405 := "1";
    null;
    r5406 := (r5405);
    r5407 := "0";
    null;
    r5408 := (r5407);
    r5409 := "1";
    null;
    r5410 := (r5409);
    r5411 := "1";
    null;
    r5412 := (r5411);
    r5413 := "0";
    null;
    r5414 := (r5413);
    r5415 := "1";
    null;
    r5416 := (r5415);
    r5417 := "1";
    null;
    r5418 := (r5417);
    r5419 := "1";
    null;
    r5420 := (r5419);
    r5421 := "0";
    null;
    r5422 := (r5421);
    r5423 := "0";
    null;
    r5424 := (r5423);
    r5425 := "1";
    null;
    r5426 := (r5425);
    r5427 := "1";
    null;
    r5428 := (r5427);
    r5429 := "1";
    null;
    r5430 := (r5429);
    r5431 := "0";
    null;
    r5432 := (r5431);
    r5433 := "0";
    null;
    r5434 := (r5433);
    r5435 := "1";
    null;
    r5436 := (r5435);
    r5437 := "1";
    null;
    r5438 := (r5437);
    r5439 := "0";
    null;
    r5440 := (r5439);
    r5441 := "0";
    null;
    r5442 := (r5441);
    r5443 := "1";
    null;
    r5444 := (r5443);
    r5445 := "0";
    null;
    r5446 := (r5445);
    r5447 := "1";
    null;
    r5448 := (r5447);
    r5449 := "0";
    null;
    r5450 := (r5449);
    r5451 := "0";
    null;
    r5452 := (r5451);
    r5453 := "1";
    null;
    r5454 := (r5453);
    r5455 := "0";
    null;
    r5456 := (r5455);
    r5457 := "0";
    null;
    r5458 := (r5457);
    r5459 := "1";
    null;
    r5460 := (r5459);
    r5461 := "1";
    null;
    r5462 := (r5461);
    r5463 := "1";
    null;
    r5464 := (r5463);
    r5465 := "1";
    null;
    r5466 := (r5465);
    r5402 := (r5404 & r5406 & r5408 & r5410 & r5412 & r5414 & r5416 & r5418 & r5420 & r5422 & r5424 & r5426 & r5428 & r5430 & r5432 & r5434 & r5436 & r5438 & r5440 & r5442 & r5444 & r5446 & r5448 & r5450 & r5452 & r5454 & r5456 & r5458 & r5460 & r5462 & r5464 & r5466);
    return r5402;
  end rewire_MetaprogrammingRW.w5b9cca4f_5401;
  function rewire_MetaprogrammingRW.w4ed8aa4a_5332 return std_logic_vector
  is
    variable r5397 : std_logic_vector(0 to 0) := (others => '0');
    variable r5396 : std_logic_vector(0 to 0) := (others => '0');
    variable r5395 : std_logic_vector(0 to 0) := (others => '0');
    variable r5394 : std_logic_vector(0 to 0) := (others => '0');
    variable r5393 : std_logic_vector(0 to 0) := (others => '0');
    variable r5392 : std_logic_vector(0 to 0) := (others => '0');
    variable r5391 : std_logic_vector(0 to 0) := (others => '0');
    variable r5390 : std_logic_vector(0 to 0) := (others => '0');
    variable r5389 : std_logic_vector(0 to 0) := (others => '0');
    variable r5388 : std_logic_vector(0 to 0) := (others => '0');
    variable r5387 : std_logic_vector(0 to 0) := (others => '0');
    variable r5386 : std_logic_vector(0 to 0) := (others => '0');
    variable r5385 : std_logic_vector(0 to 0) := (others => '0');
    variable r5384 : std_logic_vector(0 to 0) := (others => '0');
    variable r5383 : std_logic_vector(0 to 0) := (others => '0');
    variable r5382 : std_logic_vector(0 to 0) := (others => '0');
    variable r5381 : std_logic_vector(0 to 0) := (others => '0');
    variable r5380 : std_logic_vector(0 to 0) := (others => '0');
    variable r5379 : std_logic_vector(0 to 0) := (others => '0');
    variable r5378 : std_logic_vector(0 to 0) := (others => '0');
    variable r5377 : std_logic_vector(0 to 0) := (others => '0');
    variable r5376 : std_logic_vector(0 to 0) := (others => '0');
    variable r5375 : std_logic_vector(0 to 0) := (others => '0');
    variable r5374 : std_logic_vector(0 to 0) := (others => '0');
    variable r5373 : std_logic_vector(0 to 0) := (others => '0');
    variable r5372 : std_logic_vector(0 to 0) := (others => '0');
    variable r5371 : std_logic_vector(0 to 0) := (others => '0');
    variable r5370 : std_logic_vector(0 to 0) := (others => '0');
    variable r5369 : std_logic_vector(0 to 0) := (others => '0');
    variable r5368 : std_logic_vector(0 to 0) := (others => '0');
    variable r5367 : std_logic_vector(0 to 0) := (others => '0');
    variable r5366 : std_logic_vector(0 to 0) := (others => '0');
    variable r5365 : std_logic_vector(0 to 0) := (others => '0');
    variable r5364 : std_logic_vector(0 to 0) := (others => '0');
    variable r5363 : std_logic_vector(0 to 0) := (others => '0');
    variable r5362 : std_logic_vector(0 to 0) := (others => '0');
    variable r5361 : std_logic_vector(0 to 0) := (others => '0');
    variable r5360 : std_logic_vector(0 to 0) := (others => '0');
    variable r5359 : std_logic_vector(0 to 0) := (others => '0');
    variable r5358 : std_logic_vector(0 to 0) := (others => '0');
    variable r5357 : std_logic_vector(0 to 0) := (others => '0');
    variable r5356 : std_logic_vector(0 to 0) := (others => '0');
    variable r5355 : std_logic_vector(0 to 0) := (others => '0');
    variable r5354 : std_logic_vector(0 to 0) := (others => '0');
    variable r5353 : std_logic_vector(0 to 0) := (others => '0');
    variable r5352 : std_logic_vector(0 to 0) := (others => '0');
    variable r5351 : std_logic_vector(0 to 0) := (others => '0');
    variable r5350 : std_logic_vector(0 to 0) := (others => '0');
    variable r5349 : std_logic_vector(0 to 0) := (others => '0');
    variable r5348 : std_logic_vector(0 to 0) := (others => '0');
    variable r5347 : std_logic_vector(0 to 0) := (others => '0');
    variable r5346 : std_logic_vector(0 to 0) := (others => '0');
    variable r5345 : std_logic_vector(0 to 0) := (others => '0');
    variable r5344 : std_logic_vector(0 to 0) := (others => '0');
    variable r5343 : std_logic_vector(0 to 0) := (others => '0');
    variable r5342 : std_logic_vector(0 to 0) := (others => '0');
    variable r5341 : std_logic_vector(0 to 0) := (others => '0');
    variable r5340 : std_logic_vector(0 to 0) := (others => '0');
    variable r5339 : std_logic_vector(0 to 0) := (others => '0');
    variable r5338 : std_logic_vector(0 to 0) := (others => '0');
    variable r5337 : std_logic_vector(0 to 0) := (others => '0');
    variable r5336 : std_logic_vector(0 to 0) := (others => '0');
    variable r5335 : std_logic_vector(0 to 0) := (others => '0');
    variable r5334 : std_logic_vector(0 to 0) := (others => '0');
    variable r5333 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r5334 := "0";
    null;
    r5335 := (r5334);
    r5336 := "1";
    null;
    r5337 := (r5336);
    r5338 := "0";
    null;
    r5339 := (r5338);
    r5340 := "0";
    null;
    r5341 := (r5340);
    r5342 := "1";
    null;
    r5343 := (r5342);
    r5344 := "1";
    null;
    r5345 := (r5344);
    r5346 := "1";
    null;
    r5347 := (r5346);
    r5348 := "0";
    null;
    r5349 := (r5348);
    r5350 := "1";
    null;
    r5351 := (r5350);
    r5352 := "1";
    null;
    r5353 := (r5352);
    r5354 := "0";
    null;
    r5355 := (r5354);
    r5356 := "1";
    null;
    r5357 := (r5356);
    r5358 := "1";
    null;
    r5359 := (r5358);
    r5360 := "0";
    null;
    r5361 := (r5360);
    r5362 := "0";
    null;
    r5363 := (r5362);
    r5364 := "0";
    null;
    r5365 := (r5364);
    r5366 := "1";
    null;
    r5367 := (r5366);
    r5368 := "0";
    null;
    r5369 := (r5368);
    r5370 := "1";
    null;
    r5371 := (r5370);
    r5372 := "0";
    null;
    r5373 := (r5372);
    r5374 := "1";
    null;
    r5375 := (r5374);
    r5376 := "0";
    null;
    r5377 := (r5376);
    r5378 := "1";
    null;
    r5379 := (r5378);
    r5380 := "0";
    null;
    r5381 := (r5380);
    r5382 := "0";
    null;
    r5383 := (r5382);
    r5384 := "1";
    null;
    r5385 := (r5384);
    r5386 := "0";
    null;
    r5387 := (r5386);
    r5388 := "0";
    null;
    r5389 := (r5388);
    r5390 := "1";
    null;
    r5391 := (r5390);
    r5392 := "0";
    null;
    r5393 := (r5392);
    r5394 := "1";
    null;
    r5395 := (r5394);
    r5396 := "0";
    null;
    r5397 := (r5396);
    r5333 := (r5335 & r5337 & r5339 & r5341 & r5343 & r5345 & r5347 & r5349 & r5351 & r5353 & r5355 & r5357 & r5359 & r5361 & r5363 & r5365 & r5367 & r5369 & r5371 & r5373 & r5375 & r5377 & r5379 & r5381 & r5383 & r5385 & r5387 & r5389 & r5391 & r5393 & r5395 & r5397);
    return r5333;
  end rewire_MetaprogrammingRW.w4ed8aa4a_5332;
  function rewire_MetaprogrammingRW.w391c0cb3_5263 return std_logic_vector
  is
    variable r5328 : std_logic_vector(0 to 0) := (others => '0');
    variable r5327 : std_logic_vector(0 to 0) := (others => '0');
    variable r5326 : std_logic_vector(0 to 0) := (others => '0');
    variable r5325 : std_logic_vector(0 to 0) := (others => '0');
    variable r5324 : std_logic_vector(0 to 0) := (others => '0');
    variable r5323 : std_logic_vector(0 to 0) := (others => '0');
    variable r5322 : std_logic_vector(0 to 0) := (others => '0');
    variable r5321 : std_logic_vector(0 to 0) := (others => '0');
    variable r5320 : std_logic_vector(0 to 0) := (others => '0');
    variable r5319 : std_logic_vector(0 to 0) := (others => '0');
    variable r5318 : std_logic_vector(0 to 0) := (others => '0');
    variable r5317 : std_logic_vector(0 to 0) := (others => '0');
    variable r5316 : std_logic_vector(0 to 0) := (others => '0');
    variable r5315 : std_logic_vector(0 to 0) := (others => '0');
    variable r5314 : std_logic_vector(0 to 0) := (others => '0');
    variable r5313 : std_logic_vector(0 to 0) := (others => '0');
    variable r5312 : std_logic_vector(0 to 0) := (others => '0');
    variable r5311 : std_logic_vector(0 to 0) := (others => '0');
    variable r5310 : std_logic_vector(0 to 0) := (others => '0');
    variable r5309 : std_logic_vector(0 to 0) := (others => '0');
    variable r5308 : std_logic_vector(0 to 0) := (others => '0');
    variable r5307 : std_logic_vector(0 to 0) := (others => '0');
    variable r5306 : std_logic_vector(0 to 0) := (others => '0');
    variable r5305 : std_logic_vector(0 to 0) := (others => '0');
    variable r5304 : std_logic_vector(0 to 0) := (others => '0');
    variable r5303 : std_logic_vector(0 to 0) := (others => '0');
    variable r5302 : std_logic_vector(0 to 0) := (others => '0');
    variable r5301 : std_logic_vector(0 to 0) := (others => '0');
    variable r5300 : std_logic_vector(0 to 0) := (others => '0');
    variable r5299 : std_logic_vector(0 to 0) := (others => '0');
    variable r5298 : std_logic_vector(0 to 0) := (others => '0');
    variable r5297 : std_logic_vector(0 to 0) := (others => '0');
    variable r5296 : std_logic_vector(0 to 0) := (others => '0');
    variable r5295 : std_logic_vector(0 to 0) := (others => '0');
    variable r5294 : std_logic_vector(0 to 0) := (others => '0');
    variable r5293 : std_logic_vector(0 to 0) := (others => '0');
    variable r5292 : std_logic_vector(0 to 0) := (others => '0');
    variable r5291 : std_logic_vector(0 to 0) := (others => '0');
    variable r5290 : std_logic_vector(0 to 0) := (others => '0');
    variable r5289 : std_logic_vector(0 to 0) := (others => '0');
    variable r5288 : std_logic_vector(0 to 0) := (others => '0');
    variable r5287 : std_logic_vector(0 to 0) := (others => '0');
    variable r5286 : std_logic_vector(0 to 0) := (others => '0');
    variable r5285 : std_logic_vector(0 to 0) := (others => '0');
    variable r5284 : std_logic_vector(0 to 0) := (others => '0');
    variable r5283 : std_logic_vector(0 to 0) := (others => '0');
    variable r5282 : std_logic_vector(0 to 0) := (others => '0');
    variable r5281 : std_logic_vector(0 to 0) := (others => '0');
    variable r5280 : std_logic_vector(0 to 0) := (others => '0');
    variable r5279 : std_logic_vector(0 to 0) := (others => '0');
    variable r5278 : std_logic_vector(0 to 0) := (others => '0');
    variable r5277 : std_logic_vector(0 to 0) := (others => '0');
    variable r5276 : std_logic_vector(0 to 0) := (others => '0');
    variable r5275 : std_logic_vector(0 to 0) := (others => '0');
    variable r5274 : std_logic_vector(0 to 0) := (others => '0');
    variable r5273 : std_logic_vector(0 to 0) := (others => '0');
    variable r5272 : std_logic_vector(0 to 0) := (others => '0');
    variable r5271 : std_logic_vector(0 to 0) := (others => '0');
    variable r5270 : std_logic_vector(0 to 0) := (others => '0');
    variable r5269 : std_logic_vector(0 to 0) := (others => '0');
    variable r5268 : std_logic_vector(0 to 0) := (others => '0');
    variable r5267 : std_logic_vector(0 to 0) := (others => '0');
    variable r5266 : std_logic_vector(0 to 0) := (others => '0');
    variable r5265 : std_logic_vector(0 to 0) := (others => '0');
    variable r5264 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r5265 := "0";
    null;
    r5266 := (r5265);
    r5267 := "0";
    null;
    r5268 := (r5267);
    r5269 := "1";
    null;
    r5270 := (r5269);
    r5271 := "1";
    null;
    r5272 := (r5271);
    r5273 := "1";
    null;
    r5274 := (r5273);
    r5275 := "0";
    null;
    r5276 := (r5275);
    r5277 := "0";
    null;
    r5278 := (r5277);
    r5279 := "1";
    null;
    r5280 := (r5279);
    r5281 := "0";
    null;
    r5282 := (r5281);
    r5283 := "0";
    null;
    r5284 := (r5283);
    r5285 := "0";
    null;
    r5286 := (r5285);
    r5287 := "1";
    null;
    r5288 := (r5287);
    r5289 := "1";
    null;
    r5290 := (r5289);
    r5291 := "1";
    null;
    r5292 := (r5291);
    r5293 := "0";
    null;
    r5294 := (r5293);
    r5295 := "0";
    null;
    r5296 := (r5295);
    r5297 := "0";
    null;
    r5298 := (r5297);
    r5299 := "0";
    null;
    r5300 := (r5299);
    r5301 := "0";
    null;
    r5302 := (r5301);
    r5303 := "0";
    null;
    r5304 := (r5303);
    r5305 := "1";
    null;
    r5306 := (r5305);
    r5307 := "1";
    null;
    r5308 := (r5307);
    r5309 := "0";
    null;
    r5310 := (r5309);
    r5311 := "0";
    null;
    r5312 := (r5311);
    r5313 := "1";
    null;
    r5314 := (r5313);
    r5315 := "0";
    null;
    r5316 := (r5315);
    r5317 := "1";
    null;
    r5318 := (r5317);
    r5319 := "1";
    null;
    r5320 := (r5319);
    r5321 := "0";
    null;
    r5322 := (r5321);
    r5323 := "0";
    null;
    r5324 := (r5323);
    r5325 := "1";
    null;
    r5326 := (r5325);
    r5327 := "1";
    null;
    r5328 := (r5327);
    r5264 := (r5266 & r5268 & r5270 & r5272 & r5274 & r5276 & r5278 & r5280 & r5282 & r5284 & r5286 & r5288 & r5290 & r5292 & r5294 & r5296 & r5298 & r5300 & r5302 & r5304 & r5306 & r5308 & r5310 & r5312 & r5314 & r5316 & r5318 & r5320 & r5322 & r5324 & r5326 & r5328);
    return r5264;
  end rewire_MetaprogrammingRW.w391c0cb3_5263;
  function rewire_MetaprogrammingRW.w34b0bcb5_5194 return std_logic_vector
  is
    variable r5259 : std_logic_vector(0 to 0) := (others => '0');
    variable r5258 : std_logic_vector(0 to 0) := (others => '0');
    variable r5257 : std_logic_vector(0 to 0) := (others => '0');
    variable r5256 : std_logic_vector(0 to 0) := (others => '0');
    variable r5255 : std_logic_vector(0 to 0) := (others => '0');
    variable r5254 : std_logic_vector(0 to 0) := (others => '0');
    variable r5253 : std_logic_vector(0 to 0) := (others => '0');
    variable r5252 : std_logic_vector(0 to 0) := (others => '0');
    variable r5251 : std_logic_vector(0 to 0) := (others => '0');
    variable r5250 : std_logic_vector(0 to 0) := (others => '0');
    variable r5249 : std_logic_vector(0 to 0) := (others => '0');
    variable r5248 : std_logic_vector(0 to 0) := (others => '0');
    variable r5247 : std_logic_vector(0 to 0) := (others => '0');
    variable r5246 : std_logic_vector(0 to 0) := (others => '0');
    variable r5245 : std_logic_vector(0 to 0) := (others => '0');
    variable r5244 : std_logic_vector(0 to 0) := (others => '0');
    variable r5243 : std_logic_vector(0 to 0) := (others => '0');
    variable r5242 : std_logic_vector(0 to 0) := (others => '0');
    variable r5241 : std_logic_vector(0 to 0) := (others => '0');
    variable r5240 : std_logic_vector(0 to 0) := (others => '0');
    variable r5239 : std_logic_vector(0 to 0) := (others => '0');
    variable r5238 : std_logic_vector(0 to 0) := (others => '0');
    variable r5237 : std_logic_vector(0 to 0) := (others => '0');
    variable r5236 : std_logic_vector(0 to 0) := (others => '0');
    variable r5235 : std_logic_vector(0 to 0) := (others => '0');
    variable r5234 : std_logic_vector(0 to 0) := (others => '0');
    variable r5233 : std_logic_vector(0 to 0) := (others => '0');
    variable r5232 : std_logic_vector(0 to 0) := (others => '0');
    variable r5231 : std_logic_vector(0 to 0) := (others => '0');
    variable r5230 : std_logic_vector(0 to 0) := (others => '0');
    variable r5229 : std_logic_vector(0 to 0) := (others => '0');
    variable r5228 : std_logic_vector(0 to 0) := (others => '0');
    variable r5227 : std_logic_vector(0 to 0) := (others => '0');
    variable r5226 : std_logic_vector(0 to 0) := (others => '0');
    variable r5225 : std_logic_vector(0 to 0) := (others => '0');
    variable r5224 : std_logic_vector(0 to 0) := (others => '0');
    variable r5223 : std_logic_vector(0 to 0) := (others => '0');
    variable r5222 : std_logic_vector(0 to 0) := (others => '0');
    variable r5221 : std_logic_vector(0 to 0) := (others => '0');
    variable r5220 : std_logic_vector(0 to 0) := (others => '0');
    variable r5219 : std_logic_vector(0 to 0) := (others => '0');
    variable r5218 : std_logic_vector(0 to 0) := (others => '0');
    variable r5217 : std_logic_vector(0 to 0) := (others => '0');
    variable r5216 : std_logic_vector(0 to 0) := (others => '0');
    variable r5215 : std_logic_vector(0 to 0) := (others => '0');
    variable r5214 : std_logic_vector(0 to 0) := (others => '0');
    variable r5213 : std_logic_vector(0 to 0) := (others => '0');
    variable r5212 : std_logic_vector(0 to 0) := (others => '0');
    variable r5211 : std_logic_vector(0 to 0) := (others => '0');
    variable r5210 : std_logic_vector(0 to 0) := (others => '0');
    variable r5209 : std_logic_vector(0 to 0) := (others => '0');
    variable r5208 : std_logic_vector(0 to 0) := (others => '0');
    variable r5207 : std_logic_vector(0 to 0) := (others => '0');
    variable r5206 : std_logic_vector(0 to 0) := (others => '0');
    variable r5205 : std_logic_vector(0 to 0) := (others => '0');
    variable r5204 : std_logic_vector(0 to 0) := (others => '0');
    variable r5203 : std_logic_vector(0 to 0) := (others => '0');
    variable r5202 : std_logic_vector(0 to 0) := (others => '0');
    variable r5201 : std_logic_vector(0 to 0) := (others => '0');
    variable r5200 : std_logic_vector(0 to 0) := (others => '0');
    variable r5199 : std_logic_vector(0 to 0) := (others => '0');
    variable r5198 : std_logic_vector(0 to 0) := (others => '0');
    variable r5197 : std_logic_vector(0 to 0) := (others => '0');
    variable r5196 : std_logic_vector(0 to 0) := (others => '0');
    variable r5195 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r5196 := "0";
    null;
    r5197 := (r5196);
    r5198 := "0";
    null;
    r5199 := (r5198);
    r5200 := "1";
    null;
    r5201 := (r5200);
    r5202 := "1";
    null;
    r5203 := (r5202);
    r5204 := "0";
    null;
    r5205 := (r5204);
    r5206 := "1";
    null;
    r5207 := (r5206);
    r5208 := "0";
    null;
    r5209 := (r5208);
    r5210 := "0";
    null;
    r5211 := (r5210);
    r5212 := "1";
    null;
    r5213 := (r5212);
    r5214 := "0";
    null;
    r5215 := (r5214);
    r5216 := "1";
    null;
    r5217 := (r5216);
    r5218 := "1";
    null;
    r5219 := (r5218);
    r5220 := "0";
    null;
    r5221 := (r5220);
    r5222 := "0";
    null;
    r5223 := (r5222);
    r5224 := "0";
    null;
    r5225 := (r5224);
    r5226 := "0";
    null;
    r5227 := (r5226);
    r5228 := "1";
    null;
    r5229 := (r5228);
    r5230 := "0";
    null;
    r5231 := (r5230);
    r5232 := "1";
    null;
    r5233 := (r5232);
    r5234 := "1";
    null;
    r5235 := (r5234);
    r5236 := "1";
    null;
    r5237 := (r5236);
    r5238 := "1";
    null;
    r5239 := (r5238);
    r5240 := "0";
    null;
    r5241 := (r5240);
    r5242 := "0";
    null;
    r5243 := (r5242);
    r5244 := "1";
    null;
    r5245 := (r5244);
    r5246 := "0";
    null;
    r5247 := (r5246);
    r5248 := "1";
    null;
    r5249 := (r5248);
    r5250 := "1";
    null;
    r5251 := (r5250);
    r5252 := "0";
    null;
    r5253 := (r5252);
    r5254 := "1";
    null;
    r5255 := (r5254);
    r5256 := "0";
    null;
    r5257 := (r5256);
    r5258 := "1";
    null;
    r5259 := (r5258);
    r5195 := (r5197 & r5199 & r5201 & r5203 & r5205 & r5207 & r5209 & r5211 & r5213 & r5215 & r5217 & r5219 & r5221 & r5223 & r5225 & r5227 & r5229 & r5231 & r5233 & r5235 & r5237 & r5239 & r5241 & r5243 & r5245 & r5247 & r5249 & r5251 & r5253 & r5255 & r5257 & r5259);
    return r5195;
  end rewire_MetaprogrammingRW.w34b0bcb5_5194;
  function rewire_MetaprogrammingRW.w2748774c_5125 return std_logic_vector
  is
    variable r5190 : std_logic_vector(0 to 0) := (others => '0');
    variable r5189 : std_logic_vector(0 to 0) := (others => '0');
    variable r5188 : std_logic_vector(0 to 0) := (others => '0');
    variable r5187 : std_logic_vector(0 to 0) := (others => '0');
    variable r5186 : std_logic_vector(0 to 0) := (others => '0');
    variable r5185 : std_logic_vector(0 to 0) := (others => '0');
    variable r5184 : std_logic_vector(0 to 0) := (others => '0');
    variable r5183 : std_logic_vector(0 to 0) := (others => '0');
    variable r5182 : std_logic_vector(0 to 0) := (others => '0');
    variable r5181 : std_logic_vector(0 to 0) := (others => '0');
    variable r5180 : std_logic_vector(0 to 0) := (others => '0');
    variable r5179 : std_logic_vector(0 to 0) := (others => '0');
    variable r5178 : std_logic_vector(0 to 0) := (others => '0');
    variable r5177 : std_logic_vector(0 to 0) := (others => '0');
    variable r5176 : std_logic_vector(0 to 0) := (others => '0');
    variable r5175 : std_logic_vector(0 to 0) := (others => '0');
    variable r5174 : std_logic_vector(0 to 0) := (others => '0');
    variable r5173 : std_logic_vector(0 to 0) := (others => '0');
    variable r5172 : std_logic_vector(0 to 0) := (others => '0');
    variable r5171 : std_logic_vector(0 to 0) := (others => '0');
    variable r5170 : std_logic_vector(0 to 0) := (others => '0');
    variable r5169 : std_logic_vector(0 to 0) := (others => '0');
    variable r5168 : std_logic_vector(0 to 0) := (others => '0');
    variable r5167 : std_logic_vector(0 to 0) := (others => '0');
    variable r5166 : std_logic_vector(0 to 0) := (others => '0');
    variable r5165 : std_logic_vector(0 to 0) := (others => '0');
    variable r5164 : std_logic_vector(0 to 0) := (others => '0');
    variable r5163 : std_logic_vector(0 to 0) := (others => '0');
    variable r5162 : std_logic_vector(0 to 0) := (others => '0');
    variable r5161 : std_logic_vector(0 to 0) := (others => '0');
    variable r5160 : std_logic_vector(0 to 0) := (others => '0');
    variable r5159 : std_logic_vector(0 to 0) := (others => '0');
    variable r5158 : std_logic_vector(0 to 0) := (others => '0');
    variable r5157 : std_logic_vector(0 to 0) := (others => '0');
    variable r5156 : std_logic_vector(0 to 0) := (others => '0');
    variable r5155 : std_logic_vector(0 to 0) := (others => '0');
    variable r5154 : std_logic_vector(0 to 0) := (others => '0');
    variable r5153 : std_logic_vector(0 to 0) := (others => '0');
    variable r5152 : std_logic_vector(0 to 0) := (others => '0');
    variable r5151 : std_logic_vector(0 to 0) := (others => '0');
    variable r5150 : std_logic_vector(0 to 0) := (others => '0');
    variable r5149 : std_logic_vector(0 to 0) := (others => '0');
    variable r5148 : std_logic_vector(0 to 0) := (others => '0');
    variable r5147 : std_logic_vector(0 to 0) := (others => '0');
    variable r5146 : std_logic_vector(0 to 0) := (others => '0');
    variable r5145 : std_logic_vector(0 to 0) := (others => '0');
    variable r5144 : std_logic_vector(0 to 0) := (others => '0');
    variable r5143 : std_logic_vector(0 to 0) := (others => '0');
    variable r5142 : std_logic_vector(0 to 0) := (others => '0');
    variable r5141 : std_logic_vector(0 to 0) := (others => '0');
    variable r5140 : std_logic_vector(0 to 0) := (others => '0');
    variable r5139 : std_logic_vector(0 to 0) := (others => '0');
    variable r5138 : std_logic_vector(0 to 0) := (others => '0');
    variable r5137 : std_logic_vector(0 to 0) := (others => '0');
    variable r5136 : std_logic_vector(0 to 0) := (others => '0');
    variable r5135 : std_logic_vector(0 to 0) := (others => '0');
    variable r5134 : std_logic_vector(0 to 0) := (others => '0');
    variable r5133 : std_logic_vector(0 to 0) := (others => '0');
    variable r5132 : std_logic_vector(0 to 0) := (others => '0');
    variable r5131 : std_logic_vector(0 to 0) := (others => '0');
    variable r5130 : std_logic_vector(0 to 0) := (others => '0');
    variable r5129 : std_logic_vector(0 to 0) := (others => '0');
    variable r5128 : std_logic_vector(0 to 0) := (others => '0');
    variable r5127 : std_logic_vector(0 to 0) := (others => '0');
    variable r5126 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r5127 := "0";
    null;
    r5128 := (r5127);
    r5129 := "0";
    null;
    r5130 := (r5129);
    r5131 := "1";
    null;
    r5132 := (r5131);
    r5133 := "0";
    null;
    r5134 := (r5133);
    r5135 := "0";
    null;
    r5136 := (r5135);
    r5137 := "1";
    null;
    r5138 := (r5137);
    r5139 := "1";
    null;
    r5140 := (r5139);
    r5141 := "1";
    null;
    r5142 := (r5141);
    r5143 := "0";
    null;
    r5144 := (r5143);
    r5145 := "1";
    null;
    r5146 := (r5145);
    r5147 := "0";
    null;
    r5148 := (r5147);
    r5149 := "0";
    null;
    r5150 := (r5149);
    r5151 := "1";
    null;
    r5152 := (r5151);
    r5153 := "0";
    null;
    r5154 := (r5153);
    r5155 := "0";
    null;
    r5156 := (r5155);
    r5157 := "0";
    null;
    r5158 := (r5157);
    r5159 := "0";
    null;
    r5160 := (r5159);
    r5161 := "1";
    null;
    r5162 := (r5161);
    r5163 := "1";
    null;
    r5164 := (r5163);
    r5165 := "1";
    null;
    r5166 := (r5165);
    r5167 := "0";
    null;
    r5168 := (r5167);
    r5169 := "1";
    null;
    r5170 := (r5169);
    r5171 := "1";
    null;
    r5172 := (r5171);
    r5173 := "1";
    null;
    r5174 := (r5173);
    r5175 := "0";
    null;
    r5176 := (r5175);
    r5177 := "1";
    null;
    r5178 := (r5177);
    r5179 := "0";
    null;
    r5180 := (r5179);
    r5181 := "0";
    null;
    r5182 := (r5181);
    r5183 := "1";
    null;
    r5184 := (r5183);
    r5185 := "1";
    null;
    r5186 := (r5185);
    r5187 := "0";
    null;
    r5188 := (r5187);
    r5189 := "0";
    null;
    r5190 := (r5189);
    r5126 := (r5128 & r5130 & r5132 & r5134 & r5136 & r5138 & r5140 & r5142 & r5144 & r5146 & r5148 & r5150 & r5152 & r5154 & r5156 & r5158 & r5160 & r5162 & r5164 & r5166 & r5168 & r5170 & r5172 & r5174 & r5176 & r5178 & r5180 & r5182 & r5184 & r5186 & r5188 & r5190);
    return r5126;
  end rewire_MetaprogrammingRW.w2748774c_5125;
  function rewire_MetaprogrammingRW.w1e376c08_5056 return std_logic_vector
  is
    variable r5121 : std_logic_vector(0 to 0) := (others => '0');
    variable r5120 : std_logic_vector(0 to 0) := (others => '0');
    variable r5119 : std_logic_vector(0 to 0) := (others => '0');
    variable r5118 : std_logic_vector(0 to 0) := (others => '0');
    variable r5117 : std_logic_vector(0 to 0) := (others => '0');
    variable r5116 : std_logic_vector(0 to 0) := (others => '0');
    variable r5115 : std_logic_vector(0 to 0) := (others => '0');
    variable r5114 : std_logic_vector(0 to 0) := (others => '0');
    variable r5113 : std_logic_vector(0 to 0) := (others => '0');
    variable r5112 : std_logic_vector(0 to 0) := (others => '0');
    variable r5111 : std_logic_vector(0 to 0) := (others => '0');
    variable r5110 : std_logic_vector(0 to 0) := (others => '0');
    variable r5109 : std_logic_vector(0 to 0) := (others => '0');
    variable r5108 : std_logic_vector(0 to 0) := (others => '0');
    variable r5107 : std_logic_vector(0 to 0) := (others => '0');
    variable r5106 : std_logic_vector(0 to 0) := (others => '0');
    variable r5105 : std_logic_vector(0 to 0) := (others => '0');
    variable r5104 : std_logic_vector(0 to 0) := (others => '0');
    variable r5103 : std_logic_vector(0 to 0) := (others => '0');
    variable r5102 : std_logic_vector(0 to 0) := (others => '0');
    variable r5101 : std_logic_vector(0 to 0) := (others => '0');
    variable r5100 : std_logic_vector(0 to 0) := (others => '0');
    variable r5099 : std_logic_vector(0 to 0) := (others => '0');
    variable r5098 : std_logic_vector(0 to 0) := (others => '0');
    variable r5097 : std_logic_vector(0 to 0) := (others => '0');
    variable r5096 : std_logic_vector(0 to 0) := (others => '0');
    variable r5095 : std_logic_vector(0 to 0) := (others => '0');
    variable r5094 : std_logic_vector(0 to 0) := (others => '0');
    variable r5093 : std_logic_vector(0 to 0) := (others => '0');
    variable r5092 : std_logic_vector(0 to 0) := (others => '0');
    variable r5091 : std_logic_vector(0 to 0) := (others => '0');
    variable r5090 : std_logic_vector(0 to 0) := (others => '0');
    variable r5089 : std_logic_vector(0 to 0) := (others => '0');
    variable r5088 : std_logic_vector(0 to 0) := (others => '0');
    variable r5087 : std_logic_vector(0 to 0) := (others => '0');
    variable r5086 : std_logic_vector(0 to 0) := (others => '0');
    variable r5085 : std_logic_vector(0 to 0) := (others => '0');
    variable r5084 : std_logic_vector(0 to 0) := (others => '0');
    variable r5083 : std_logic_vector(0 to 0) := (others => '0');
    variable r5082 : std_logic_vector(0 to 0) := (others => '0');
    variable r5081 : std_logic_vector(0 to 0) := (others => '0');
    variable r5080 : std_logic_vector(0 to 0) := (others => '0');
    variable r5079 : std_logic_vector(0 to 0) := (others => '0');
    variable r5078 : std_logic_vector(0 to 0) := (others => '0');
    variable r5077 : std_logic_vector(0 to 0) := (others => '0');
    variable r5076 : std_logic_vector(0 to 0) := (others => '0');
    variable r5075 : std_logic_vector(0 to 0) := (others => '0');
    variable r5074 : std_logic_vector(0 to 0) := (others => '0');
    variable r5073 : std_logic_vector(0 to 0) := (others => '0');
    variable r5072 : std_logic_vector(0 to 0) := (others => '0');
    variable r5071 : std_logic_vector(0 to 0) := (others => '0');
    variable r5070 : std_logic_vector(0 to 0) := (others => '0');
    variable r5069 : std_logic_vector(0 to 0) := (others => '0');
    variable r5068 : std_logic_vector(0 to 0) := (others => '0');
    variable r5067 : std_logic_vector(0 to 0) := (others => '0');
    variable r5066 : std_logic_vector(0 to 0) := (others => '0');
    variable r5065 : std_logic_vector(0 to 0) := (others => '0');
    variable r5064 : std_logic_vector(0 to 0) := (others => '0');
    variable r5063 : std_logic_vector(0 to 0) := (others => '0');
    variable r5062 : std_logic_vector(0 to 0) := (others => '0');
    variable r5061 : std_logic_vector(0 to 0) := (others => '0');
    variable r5060 : std_logic_vector(0 to 0) := (others => '0');
    variable r5059 : std_logic_vector(0 to 0) := (others => '0');
    variable r5058 : std_logic_vector(0 to 0) := (others => '0');
    variable r5057 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r5058 := "0";
    null;
    r5059 := (r5058);
    r5060 := "0";
    null;
    r5061 := (r5060);
    r5062 := "0";
    null;
    r5063 := (r5062);
    r5064 := "1";
    null;
    r5065 := (r5064);
    r5066 := "1";
    null;
    r5067 := (r5066);
    r5068 := "1";
    null;
    r5069 := (r5068);
    r5070 := "1";
    null;
    r5071 := (r5070);
    r5072 := "0";
    null;
    r5073 := (r5072);
    r5074 := "0";
    null;
    r5075 := (r5074);
    r5076 := "0";
    null;
    r5077 := (r5076);
    r5078 := "1";
    null;
    r5079 := (r5078);
    r5080 := "1";
    null;
    r5081 := (r5080);
    r5082 := "0";
    null;
    r5083 := (r5082);
    r5084 := "1";
    null;
    r5085 := (r5084);
    r5086 := "1";
    null;
    r5087 := (r5086);
    r5088 := "1";
    null;
    r5089 := (r5088);
    r5090 := "0";
    null;
    r5091 := (r5090);
    r5092 := "1";
    null;
    r5093 := (r5092);
    r5094 := "1";
    null;
    r5095 := (r5094);
    r5096 := "0";
    null;
    r5097 := (r5096);
    r5098 := "1";
    null;
    r5099 := (r5098);
    r5100 := "1";
    null;
    r5101 := (r5100);
    r5102 := "0";
    null;
    r5103 := (r5102);
    r5104 := "0";
    null;
    r5105 := (r5104);
    r5106 := "0";
    null;
    r5107 := (r5106);
    r5108 := "0";
    null;
    r5109 := (r5108);
    r5110 := "0";
    null;
    r5111 := (r5110);
    r5112 := "0";
    null;
    r5113 := (r5112);
    r5114 := "1";
    null;
    r5115 := (r5114);
    r5116 := "0";
    null;
    r5117 := (r5116);
    r5118 := "0";
    null;
    r5119 := (r5118);
    r5120 := "0";
    null;
    r5121 := (r5120);
    r5057 := (r5059 & r5061 & r5063 & r5065 & r5067 & r5069 & r5071 & r5073 & r5075 & r5077 & r5079 & r5081 & r5083 & r5085 & r5087 & r5089 & r5091 & r5093 & r5095 & r5097 & r5099 & r5101 & r5103 & r5105 & r5107 & r5109 & r5111 & r5113 & r5115 & r5117 & r5119 & r5121);
    return r5057;
  end rewire_MetaprogrammingRW.w1e376c08_5056;
  function rewire_MetaprogrammingRW.w19a4c116_4987 return std_logic_vector
  is
    variable r5052 : std_logic_vector(0 to 0) := (others => '0');
    variable r5051 : std_logic_vector(0 to 0) := (others => '0');
    variable r5050 : std_logic_vector(0 to 0) := (others => '0');
    variable r5049 : std_logic_vector(0 to 0) := (others => '0');
    variable r5048 : std_logic_vector(0 to 0) := (others => '0');
    variable r5047 : std_logic_vector(0 to 0) := (others => '0');
    variable r5046 : std_logic_vector(0 to 0) := (others => '0');
    variable r5045 : std_logic_vector(0 to 0) := (others => '0');
    variable r5044 : std_logic_vector(0 to 0) := (others => '0');
    variable r5043 : std_logic_vector(0 to 0) := (others => '0');
    variable r5042 : std_logic_vector(0 to 0) := (others => '0');
    variable r5041 : std_logic_vector(0 to 0) := (others => '0');
    variable r5040 : std_logic_vector(0 to 0) := (others => '0');
    variable r5039 : std_logic_vector(0 to 0) := (others => '0');
    variable r5038 : std_logic_vector(0 to 0) := (others => '0');
    variable r5037 : std_logic_vector(0 to 0) := (others => '0');
    variable r5036 : std_logic_vector(0 to 0) := (others => '0');
    variable r5035 : std_logic_vector(0 to 0) := (others => '0');
    variable r5034 : std_logic_vector(0 to 0) := (others => '0');
    variable r5033 : std_logic_vector(0 to 0) := (others => '0');
    variable r5032 : std_logic_vector(0 to 0) := (others => '0');
    variable r5031 : std_logic_vector(0 to 0) := (others => '0');
    variable r5030 : std_logic_vector(0 to 0) := (others => '0');
    variable r5029 : std_logic_vector(0 to 0) := (others => '0');
    variable r5028 : std_logic_vector(0 to 0) := (others => '0');
    variable r5027 : std_logic_vector(0 to 0) := (others => '0');
    variable r5026 : std_logic_vector(0 to 0) := (others => '0');
    variable r5025 : std_logic_vector(0 to 0) := (others => '0');
    variable r5024 : std_logic_vector(0 to 0) := (others => '0');
    variable r5023 : std_logic_vector(0 to 0) := (others => '0');
    variable r5022 : std_logic_vector(0 to 0) := (others => '0');
    variable r5021 : std_logic_vector(0 to 0) := (others => '0');
    variable r5020 : std_logic_vector(0 to 0) := (others => '0');
    variable r5019 : std_logic_vector(0 to 0) := (others => '0');
    variable r5018 : std_logic_vector(0 to 0) := (others => '0');
    variable r5017 : std_logic_vector(0 to 0) := (others => '0');
    variable r5016 : std_logic_vector(0 to 0) := (others => '0');
    variable r5015 : std_logic_vector(0 to 0) := (others => '0');
    variable r5014 : std_logic_vector(0 to 0) := (others => '0');
    variable r5013 : std_logic_vector(0 to 0) := (others => '0');
    variable r5012 : std_logic_vector(0 to 0) := (others => '0');
    variable r5011 : std_logic_vector(0 to 0) := (others => '0');
    variable r5010 : std_logic_vector(0 to 0) := (others => '0');
    variable r5009 : std_logic_vector(0 to 0) := (others => '0');
    variable r5008 : std_logic_vector(0 to 0) := (others => '0');
    variable r5007 : std_logic_vector(0 to 0) := (others => '0');
    variable r5006 : std_logic_vector(0 to 0) := (others => '0');
    variable r5005 : std_logic_vector(0 to 0) := (others => '0');
    variable r5004 : std_logic_vector(0 to 0) := (others => '0');
    variable r5003 : std_logic_vector(0 to 0) := (others => '0');
    variable r5002 : std_logic_vector(0 to 0) := (others => '0');
    variable r5001 : std_logic_vector(0 to 0) := (others => '0');
    variable r5000 : std_logic_vector(0 to 0) := (others => '0');
    variable r4999 : std_logic_vector(0 to 0) := (others => '0');
    variable r4998 : std_logic_vector(0 to 0) := (others => '0');
    variable r4997 : std_logic_vector(0 to 0) := (others => '0');
    variable r4996 : std_logic_vector(0 to 0) := (others => '0');
    variable r4995 : std_logic_vector(0 to 0) := (others => '0');
    variable r4994 : std_logic_vector(0 to 0) := (others => '0');
    variable r4993 : std_logic_vector(0 to 0) := (others => '0');
    variable r4992 : std_logic_vector(0 to 0) := (others => '0');
    variable r4991 : std_logic_vector(0 to 0) := (others => '0');
    variable r4990 : std_logic_vector(0 to 0) := (others => '0');
    variable r4989 : std_logic_vector(0 to 0) := (others => '0');
    variable r4988 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r4989 := "0";
    null;
    r4990 := (r4989);
    r4991 := "0";
    null;
    r4992 := (r4991);
    r4993 := "0";
    null;
    r4994 := (r4993);
    r4995 := "1";
    null;
    r4996 := (r4995);
    r4997 := "1";
    null;
    r4998 := (r4997);
    r4999 := "0";
    null;
    r5000 := (r4999);
    r5001 := "0";
    null;
    r5002 := (r5001);
    r5003 := "1";
    null;
    r5004 := (r5003);
    r5005 := "1";
    null;
    r5006 := (r5005);
    r5007 := "0";
    null;
    r5008 := (r5007);
    r5009 := "1";
    null;
    r5010 := (r5009);
    r5011 := "0";
    null;
    r5012 := (r5011);
    r5013 := "0";
    null;
    r5014 := (r5013);
    r5015 := "1";
    null;
    r5016 := (r5015);
    r5017 := "0";
    null;
    r5018 := (r5017);
    r5019 := "0";
    null;
    r5020 := (r5019);
    r5021 := "1";
    null;
    r5022 := (r5021);
    r5023 := "1";
    null;
    r5024 := (r5023);
    r5025 := "0";
    null;
    r5026 := (r5025);
    r5027 := "0";
    null;
    r5028 := (r5027);
    r5029 := "0";
    null;
    r5030 := (r5029);
    r5031 := "0";
    null;
    r5032 := (r5031);
    r5033 := "0";
    null;
    r5034 := (r5033);
    r5035 := "1";
    null;
    r5036 := (r5035);
    r5037 := "0";
    null;
    r5038 := (r5037);
    r5039 := "0";
    null;
    r5040 := (r5039);
    r5041 := "0";
    null;
    r5042 := (r5041);
    r5043 := "1";
    null;
    r5044 := (r5043);
    r5045 := "0";
    null;
    r5046 := (r5045);
    r5047 := "1";
    null;
    r5048 := (r5047);
    r5049 := "1";
    null;
    r5050 := (r5049);
    r5051 := "0";
    null;
    r5052 := (r5051);
    r4988 := (r4990 & r4992 & r4994 & r4996 & r4998 & r5000 & r5002 & r5004 & r5006 & r5008 & r5010 & r5012 & r5014 & r5016 & r5018 & r5020 & r5022 & r5024 & r5026 & r5028 & r5030 & r5032 & r5034 & r5036 & r5038 & r5040 & r5042 & r5044 & r5046 & r5048 & r5050 & r5052);
    return r4988;
  end rewire_MetaprogrammingRW.w19a4c116_4987;
  function rewire_MetaprogrammingRW.w106aa070_4918 return std_logic_vector
  is
    variable r4983 : std_logic_vector(0 to 0) := (others => '0');
    variable r4982 : std_logic_vector(0 to 0) := (others => '0');
    variable r4981 : std_logic_vector(0 to 0) := (others => '0');
    variable r4980 : std_logic_vector(0 to 0) := (others => '0');
    variable r4979 : std_logic_vector(0 to 0) := (others => '0');
    variable r4978 : std_logic_vector(0 to 0) := (others => '0');
    variable r4977 : std_logic_vector(0 to 0) := (others => '0');
    variable r4976 : std_logic_vector(0 to 0) := (others => '0');
    variable r4975 : std_logic_vector(0 to 0) := (others => '0');
    variable r4974 : std_logic_vector(0 to 0) := (others => '0');
    variable r4973 : std_logic_vector(0 to 0) := (others => '0');
    variable r4972 : std_logic_vector(0 to 0) := (others => '0');
    variable r4971 : std_logic_vector(0 to 0) := (others => '0');
    variable r4970 : std_logic_vector(0 to 0) := (others => '0');
    variable r4969 : std_logic_vector(0 to 0) := (others => '0');
    variable r4968 : std_logic_vector(0 to 0) := (others => '0');
    variable r4967 : std_logic_vector(0 to 0) := (others => '0');
    variable r4966 : std_logic_vector(0 to 0) := (others => '0');
    variable r4965 : std_logic_vector(0 to 0) := (others => '0');
    variable r4964 : std_logic_vector(0 to 0) := (others => '0');
    variable r4963 : std_logic_vector(0 to 0) := (others => '0');
    variable r4962 : std_logic_vector(0 to 0) := (others => '0');
    variable r4961 : std_logic_vector(0 to 0) := (others => '0');
    variable r4960 : std_logic_vector(0 to 0) := (others => '0');
    variable r4959 : std_logic_vector(0 to 0) := (others => '0');
    variable r4958 : std_logic_vector(0 to 0) := (others => '0');
    variable r4957 : std_logic_vector(0 to 0) := (others => '0');
    variable r4956 : std_logic_vector(0 to 0) := (others => '0');
    variable r4955 : std_logic_vector(0 to 0) := (others => '0');
    variable r4954 : std_logic_vector(0 to 0) := (others => '0');
    variable r4953 : std_logic_vector(0 to 0) := (others => '0');
    variable r4952 : std_logic_vector(0 to 0) := (others => '0');
    variable r4951 : std_logic_vector(0 to 0) := (others => '0');
    variable r4950 : std_logic_vector(0 to 0) := (others => '0');
    variable r4949 : std_logic_vector(0 to 0) := (others => '0');
    variable r4948 : std_logic_vector(0 to 0) := (others => '0');
    variable r4947 : std_logic_vector(0 to 0) := (others => '0');
    variable r4946 : std_logic_vector(0 to 0) := (others => '0');
    variable r4945 : std_logic_vector(0 to 0) := (others => '0');
    variable r4944 : std_logic_vector(0 to 0) := (others => '0');
    variable r4943 : std_logic_vector(0 to 0) := (others => '0');
    variable r4942 : std_logic_vector(0 to 0) := (others => '0');
    variable r4941 : std_logic_vector(0 to 0) := (others => '0');
    variable r4940 : std_logic_vector(0 to 0) := (others => '0');
    variable r4939 : std_logic_vector(0 to 0) := (others => '0');
    variable r4938 : std_logic_vector(0 to 0) := (others => '0');
    variable r4937 : std_logic_vector(0 to 0) := (others => '0');
    variable r4936 : std_logic_vector(0 to 0) := (others => '0');
    variable r4935 : std_logic_vector(0 to 0) := (others => '0');
    variable r4934 : std_logic_vector(0 to 0) := (others => '0');
    variable r4933 : std_logic_vector(0 to 0) := (others => '0');
    variable r4932 : std_logic_vector(0 to 0) := (others => '0');
    variable r4931 : std_logic_vector(0 to 0) := (others => '0');
    variable r4930 : std_logic_vector(0 to 0) := (others => '0');
    variable r4929 : std_logic_vector(0 to 0) := (others => '0');
    variable r4928 : std_logic_vector(0 to 0) := (others => '0');
    variable r4927 : std_logic_vector(0 to 0) := (others => '0');
    variable r4926 : std_logic_vector(0 to 0) := (others => '0');
    variable r4925 : std_logic_vector(0 to 0) := (others => '0');
    variable r4924 : std_logic_vector(0 to 0) := (others => '0');
    variable r4923 : std_logic_vector(0 to 0) := (others => '0');
    variable r4922 : std_logic_vector(0 to 0) := (others => '0');
    variable r4921 : std_logic_vector(0 to 0) := (others => '0');
    variable r4920 : std_logic_vector(0 to 0) := (others => '0');
    variable r4919 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r4920 := "0";
    null;
    r4921 := (r4920);
    r4922 := "0";
    null;
    r4923 := (r4922);
    r4924 := "0";
    null;
    r4925 := (r4924);
    r4926 := "1";
    null;
    r4927 := (r4926);
    r4928 := "0";
    null;
    r4929 := (r4928);
    r4930 := "0";
    null;
    r4931 := (r4930);
    r4932 := "0";
    null;
    r4933 := (r4932);
    r4934 := "0";
    null;
    r4935 := (r4934);
    r4936 := "0";
    null;
    r4937 := (r4936);
    r4938 := "1";
    null;
    r4939 := (r4938);
    r4940 := "1";
    null;
    r4941 := (r4940);
    r4942 := "0";
    null;
    r4943 := (r4942);
    r4944 := "1";
    null;
    r4945 := (r4944);
    r4946 := "0";
    null;
    r4947 := (r4946);
    r4948 := "1";
    null;
    r4949 := (r4948);
    r4950 := "0";
    null;
    r4951 := (r4950);
    r4952 := "1";
    null;
    r4953 := (r4952);
    r4954 := "0";
    null;
    r4955 := (r4954);
    r4956 := "1";
    null;
    r4957 := (r4956);
    r4958 := "0";
    null;
    r4959 := (r4958);
    r4960 := "0";
    null;
    r4961 := (r4960);
    r4962 := "0";
    null;
    r4963 := (r4962);
    r4964 := "0";
    null;
    r4965 := (r4964);
    r4966 := "0";
    null;
    r4967 := (r4966);
    r4968 := "0";
    null;
    r4969 := (r4968);
    r4970 := "1";
    null;
    r4971 := (r4970);
    r4972 := "1";
    null;
    r4973 := (r4972);
    r4974 := "1";
    null;
    r4975 := (r4974);
    r4976 := "0";
    null;
    r4977 := (r4976);
    r4978 := "0";
    null;
    r4979 := (r4978);
    r4980 := "0";
    null;
    r4981 := (r4980);
    r4982 := "0";
    null;
    r4983 := (r4982);
    r4919 := (r4921 & r4923 & r4925 & r4927 & r4929 & r4931 & r4933 & r4935 & r4937 & r4939 & r4941 & r4943 & r4945 & r4947 & r4949 & r4951 & r4953 & r4955 & r4957 & r4959 & r4961 & r4963 & r4965 & r4967 & r4969 & r4971 & r4973 & r4975 & r4977 & r4979 & r4981 & r4983);
    return r4919;
  end rewire_MetaprogrammingRW.w106aa070_4918;
  function rewire_MetaprogrammingRW.wf40e3585_4849 return std_logic_vector
  is
    variable r4914 : std_logic_vector(0 to 0) := (others => '0');
    variable r4913 : std_logic_vector(0 to 0) := (others => '0');
    variable r4912 : std_logic_vector(0 to 0) := (others => '0');
    variable r4911 : std_logic_vector(0 to 0) := (others => '0');
    variable r4910 : std_logic_vector(0 to 0) := (others => '0');
    variable r4909 : std_logic_vector(0 to 0) := (others => '0');
    variable r4908 : std_logic_vector(0 to 0) := (others => '0');
    variable r4907 : std_logic_vector(0 to 0) := (others => '0');
    variable r4906 : std_logic_vector(0 to 0) := (others => '0');
    variable r4905 : std_logic_vector(0 to 0) := (others => '0');
    variable r4904 : std_logic_vector(0 to 0) := (others => '0');
    variable r4903 : std_logic_vector(0 to 0) := (others => '0');
    variable r4902 : std_logic_vector(0 to 0) := (others => '0');
    variable r4901 : std_logic_vector(0 to 0) := (others => '0');
    variable r4900 : std_logic_vector(0 to 0) := (others => '0');
    variable r4899 : std_logic_vector(0 to 0) := (others => '0');
    variable r4898 : std_logic_vector(0 to 0) := (others => '0');
    variable r4897 : std_logic_vector(0 to 0) := (others => '0');
    variable r4896 : std_logic_vector(0 to 0) := (others => '0');
    variable r4895 : std_logic_vector(0 to 0) := (others => '0');
    variable r4894 : std_logic_vector(0 to 0) := (others => '0');
    variable r4893 : std_logic_vector(0 to 0) := (others => '0');
    variable r4892 : std_logic_vector(0 to 0) := (others => '0');
    variable r4891 : std_logic_vector(0 to 0) := (others => '0');
    variable r4890 : std_logic_vector(0 to 0) := (others => '0');
    variable r4889 : std_logic_vector(0 to 0) := (others => '0');
    variable r4888 : std_logic_vector(0 to 0) := (others => '0');
    variable r4887 : std_logic_vector(0 to 0) := (others => '0');
    variable r4886 : std_logic_vector(0 to 0) := (others => '0');
    variable r4885 : std_logic_vector(0 to 0) := (others => '0');
    variable r4884 : std_logic_vector(0 to 0) := (others => '0');
    variable r4883 : std_logic_vector(0 to 0) := (others => '0');
    variable r4882 : std_logic_vector(0 to 0) := (others => '0');
    variable r4881 : std_logic_vector(0 to 0) := (others => '0');
    variable r4880 : std_logic_vector(0 to 0) := (others => '0');
    variable r4879 : std_logic_vector(0 to 0) := (others => '0');
    variable r4878 : std_logic_vector(0 to 0) := (others => '0');
    variable r4877 : std_logic_vector(0 to 0) := (others => '0');
    variable r4876 : std_logic_vector(0 to 0) := (others => '0');
    variable r4875 : std_logic_vector(0 to 0) := (others => '0');
    variable r4874 : std_logic_vector(0 to 0) := (others => '0');
    variable r4873 : std_logic_vector(0 to 0) := (others => '0');
    variable r4872 : std_logic_vector(0 to 0) := (others => '0');
    variable r4871 : std_logic_vector(0 to 0) := (others => '0');
    variable r4870 : std_logic_vector(0 to 0) := (others => '0');
    variable r4869 : std_logic_vector(0 to 0) := (others => '0');
    variable r4868 : std_logic_vector(0 to 0) := (others => '0');
    variable r4867 : std_logic_vector(0 to 0) := (others => '0');
    variable r4866 : std_logic_vector(0 to 0) := (others => '0');
    variable r4865 : std_logic_vector(0 to 0) := (others => '0');
    variable r4864 : std_logic_vector(0 to 0) := (others => '0');
    variable r4863 : std_logic_vector(0 to 0) := (others => '0');
    variable r4862 : std_logic_vector(0 to 0) := (others => '0');
    variable r4861 : std_logic_vector(0 to 0) := (others => '0');
    variable r4860 : std_logic_vector(0 to 0) := (others => '0');
    variable r4859 : std_logic_vector(0 to 0) := (others => '0');
    variable r4858 : std_logic_vector(0 to 0) := (others => '0');
    variable r4857 : std_logic_vector(0 to 0) := (others => '0');
    variable r4856 : std_logic_vector(0 to 0) := (others => '0');
    variable r4855 : std_logic_vector(0 to 0) := (others => '0');
    variable r4854 : std_logic_vector(0 to 0) := (others => '0');
    variable r4853 : std_logic_vector(0 to 0) := (others => '0');
    variable r4852 : std_logic_vector(0 to 0) := (others => '0');
    variable r4851 : std_logic_vector(0 to 0) := (others => '0');
    variable r4850 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r4851 := "1";
    null;
    r4852 := (r4851);
    r4853 := "1";
    null;
    r4854 := (r4853);
    r4855 := "1";
    null;
    r4856 := (r4855);
    r4857 := "1";
    null;
    r4858 := (r4857);
    r4859 := "0";
    null;
    r4860 := (r4859);
    r4861 := "1";
    null;
    r4862 := (r4861);
    r4863 := "0";
    null;
    r4864 := (r4863);
    r4865 := "0";
    null;
    r4866 := (r4865);
    r4867 := "0";
    null;
    r4868 := (r4867);
    r4869 := "0";
    null;
    r4870 := (r4869);
    r4871 := "0";
    null;
    r4872 := (r4871);
    r4873 := "0";
    null;
    r4874 := (r4873);
    r4875 := "1";
    null;
    r4876 := (r4875);
    r4877 := "1";
    null;
    r4878 := (r4877);
    r4879 := "1";
    null;
    r4880 := (r4879);
    r4881 := "0";
    null;
    r4882 := (r4881);
    r4883 := "0";
    null;
    r4884 := (r4883);
    r4885 := "0";
    null;
    r4886 := (r4885);
    r4887 := "1";
    null;
    r4888 := (r4887);
    r4889 := "1";
    null;
    r4890 := (r4889);
    r4891 := "0";
    null;
    r4892 := (r4891);
    r4893 := "1";
    null;
    r4894 := (r4893);
    r4895 := "0";
    null;
    r4896 := (r4895);
    r4897 := "1";
    null;
    r4898 := (r4897);
    r4899 := "1";
    null;
    r4900 := (r4899);
    r4901 := "0";
    null;
    r4902 := (r4901);
    r4903 := "0";
    null;
    r4904 := (r4903);
    r4905 := "0";
    null;
    r4906 := (r4905);
    r4907 := "0";
    null;
    r4908 := (r4907);
    r4909 := "1";
    null;
    r4910 := (r4909);
    r4911 := "0";
    null;
    r4912 := (r4911);
    r4913 := "1";
    null;
    r4914 := (r4913);
    r4850 := (r4852 & r4854 & r4856 & r4858 & r4860 & r4862 & r4864 & r4866 & r4868 & r4870 & r4872 & r4874 & r4876 & r4878 & r4880 & r4882 & r4884 & r4886 & r4888 & r4890 & r4892 & r4894 & r4896 & r4898 & r4900 & r4902 & r4904 & r4906 & r4908 & r4910 & r4912 & r4914);
    return r4850;
  end rewire_MetaprogrammingRW.wf40e3585_4849;
  function rewire_MetaprogrammingRW.wd6990624_4780 return std_logic_vector
  is
    variable r4845 : std_logic_vector(0 to 0) := (others => '0');
    variable r4844 : std_logic_vector(0 to 0) := (others => '0');
    variable r4843 : std_logic_vector(0 to 0) := (others => '0');
    variable r4842 : std_logic_vector(0 to 0) := (others => '0');
    variable r4841 : std_logic_vector(0 to 0) := (others => '0');
    variable r4840 : std_logic_vector(0 to 0) := (others => '0');
    variable r4839 : std_logic_vector(0 to 0) := (others => '0');
    variable r4838 : std_logic_vector(0 to 0) := (others => '0');
    variable r4837 : std_logic_vector(0 to 0) := (others => '0');
    variable r4836 : std_logic_vector(0 to 0) := (others => '0');
    variable r4835 : std_logic_vector(0 to 0) := (others => '0');
    variable r4834 : std_logic_vector(0 to 0) := (others => '0');
    variable r4833 : std_logic_vector(0 to 0) := (others => '0');
    variable r4832 : std_logic_vector(0 to 0) := (others => '0');
    variable r4831 : std_logic_vector(0 to 0) := (others => '0');
    variable r4830 : std_logic_vector(0 to 0) := (others => '0');
    variable r4829 : std_logic_vector(0 to 0) := (others => '0');
    variable r4828 : std_logic_vector(0 to 0) := (others => '0');
    variable r4827 : std_logic_vector(0 to 0) := (others => '0');
    variable r4826 : std_logic_vector(0 to 0) := (others => '0');
    variable r4825 : std_logic_vector(0 to 0) := (others => '0');
    variable r4824 : std_logic_vector(0 to 0) := (others => '0');
    variable r4823 : std_logic_vector(0 to 0) := (others => '0');
    variable r4822 : std_logic_vector(0 to 0) := (others => '0');
    variable r4821 : std_logic_vector(0 to 0) := (others => '0');
    variable r4820 : std_logic_vector(0 to 0) := (others => '0');
    variable r4819 : std_logic_vector(0 to 0) := (others => '0');
    variable r4818 : std_logic_vector(0 to 0) := (others => '0');
    variable r4817 : std_logic_vector(0 to 0) := (others => '0');
    variable r4816 : std_logic_vector(0 to 0) := (others => '0');
    variable r4815 : std_logic_vector(0 to 0) := (others => '0');
    variable r4814 : std_logic_vector(0 to 0) := (others => '0');
    variable r4813 : std_logic_vector(0 to 0) := (others => '0');
    variable r4812 : std_logic_vector(0 to 0) := (others => '0');
    variable r4811 : std_logic_vector(0 to 0) := (others => '0');
    variable r4810 : std_logic_vector(0 to 0) := (others => '0');
    variable r4809 : std_logic_vector(0 to 0) := (others => '0');
    variable r4808 : std_logic_vector(0 to 0) := (others => '0');
    variable r4807 : std_logic_vector(0 to 0) := (others => '0');
    variable r4806 : std_logic_vector(0 to 0) := (others => '0');
    variable r4805 : std_logic_vector(0 to 0) := (others => '0');
    variable r4804 : std_logic_vector(0 to 0) := (others => '0');
    variable r4803 : std_logic_vector(0 to 0) := (others => '0');
    variable r4802 : std_logic_vector(0 to 0) := (others => '0');
    variable r4801 : std_logic_vector(0 to 0) := (others => '0');
    variable r4800 : std_logic_vector(0 to 0) := (others => '0');
    variable r4799 : std_logic_vector(0 to 0) := (others => '0');
    variable r4798 : std_logic_vector(0 to 0) := (others => '0');
    variable r4797 : std_logic_vector(0 to 0) := (others => '0');
    variable r4796 : std_logic_vector(0 to 0) := (others => '0');
    variable r4795 : std_logic_vector(0 to 0) := (others => '0');
    variable r4794 : std_logic_vector(0 to 0) := (others => '0');
    variable r4793 : std_logic_vector(0 to 0) := (others => '0');
    variable r4792 : std_logic_vector(0 to 0) := (others => '0');
    variable r4791 : std_logic_vector(0 to 0) := (others => '0');
    variable r4790 : std_logic_vector(0 to 0) := (others => '0');
    variable r4789 : std_logic_vector(0 to 0) := (others => '0');
    variable r4788 : std_logic_vector(0 to 0) := (others => '0');
    variable r4787 : std_logic_vector(0 to 0) := (others => '0');
    variable r4786 : std_logic_vector(0 to 0) := (others => '0');
    variable r4785 : std_logic_vector(0 to 0) := (others => '0');
    variable r4784 : std_logic_vector(0 to 0) := (others => '0');
    variable r4783 : std_logic_vector(0 to 0) := (others => '0');
    variable r4782 : std_logic_vector(0 to 0) := (others => '0');
    variable r4781 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r4782 := "1";
    null;
    r4783 := (r4782);
    r4784 := "1";
    null;
    r4785 := (r4784);
    r4786 := "0";
    null;
    r4787 := (r4786);
    r4788 := "1";
    null;
    r4789 := (r4788);
    r4790 := "0";
    null;
    r4791 := (r4790);
    r4792 := "1";
    null;
    r4793 := (r4792);
    r4794 := "1";
    null;
    r4795 := (r4794);
    r4796 := "0";
    null;
    r4797 := (r4796);
    r4798 := "1";
    null;
    r4799 := (r4798);
    r4800 := "0";
    null;
    r4801 := (r4800);
    r4802 := "0";
    null;
    r4803 := (r4802);
    r4804 := "1";
    null;
    r4805 := (r4804);
    r4806 := "1";
    null;
    r4807 := (r4806);
    r4808 := "0";
    null;
    r4809 := (r4808);
    r4810 := "0";
    null;
    r4811 := (r4810);
    r4812 := "1";
    null;
    r4813 := (r4812);
    r4814 := "0";
    null;
    r4815 := (r4814);
    r4816 := "0";
    null;
    r4817 := (r4816);
    r4818 := "0";
    null;
    r4819 := (r4818);
    r4820 := "0";
    null;
    r4821 := (r4820);
    r4822 := "0";
    null;
    r4823 := (r4822);
    r4824 := "1";
    null;
    r4825 := (r4824);
    r4826 := "1";
    null;
    r4827 := (r4826);
    r4828 := "0";
    null;
    r4829 := (r4828);
    r4830 := "0";
    null;
    r4831 := (r4830);
    r4832 := "0";
    null;
    r4833 := (r4832);
    r4834 := "1";
    null;
    r4835 := (r4834);
    r4836 := "0";
    null;
    r4837 := (r4836);
    r4838 := "0";
    null;
    r4839 := (r4838);
    r4840 := "1";
    null;
    r4841 := (r4840);
    r4842 := "0";
    null;
    r4843 := (r4842);
    r4844 := "0";
    null;
    r4845 := (r4844);
    r4781 := (r4783 & r4785 & r4787 & r4789 & r4791 & r4793 & r4795 & r4797 & r4799 & r4801 & r4803 & r4805 & r4807 & r4809 & r4811 & r4813 & r4815 & r4817 & r4819 & r4821 & r4823 & r4825 & r4827 & r4829 & r4831 & r4833 & r4835 & r4837 & r4839 & r4841 & r4843 & r4845);
    return r4781;
  end rewire_MetaprogrammingRW.wd6990624_4780;
  function rewire_MetaprogrammingRW.wd192e819_4711 return std_logic_vector
  is
    variable r4776 : std_logic_vector(0 to 0) := (others => '0');
    variable r4775 : std_logic_vector(0 to 0) := (others => '0');
    variable r4774 : std_logic_vector(0 to 0) := (others => '0');
    variable r4773 : std_logic_vector(0 to 0) := (others => '0');
    variable r4772 : std_logic_vector(0 to 0) := (others => '0');
    variable r4771 : std_logic_vector(0 to 0) := (others => '0');
    variable r4770 : std_logic_vector(0 to 0) := (others => '0');
    variable r4769 : std_logic_vector(0 to 0) := (others => '0');
    variable r4768 : std_logic_vector(0 to 0) := (others => '0');
    variable r4767 : std_logic_vector(0 to 0) := (others => '0');
    variable r4766 : std_logic_vector(0 to 0) := (others => '0');
    variable r4765 : std_logic_vector(0 to 0) := (others => '0');
    variable r4764 : std_logic_vector(0 to 0) := (others => '0');
    variable r4763 : std_logic_vector(0 to 0) := (others => '0');
    variable r4762 : std_logic_vector(0 to 0) := (others => '0');
    variable r4761 : std_logic_vector(0 to 0) := (others => '0');
    variable r4760 : std_logic_vector(0 to 0) := (others => '0');
    variable r4759 : std_logic_vector(0 to 0) := (others => '0');
    variable r4758 : std_logic_vector(0 to 0) := (others => '0');
    variable r4757 : std_logic_vector(0 to 0) := (others => '0');
    variable r4756 : std_logic_vector(0 to 0) := (others => '0');
    variable r4755 : std_logic_vector(0 to 0) := (others => '0');
    variable r4754 : std_logic_vector(0 to 0) := (others => '0');
    variable r4753 : std_logic_vector(0 to 0) := (others => '0');
    variable r4752 : std_logic_vector(0 to 0) := (others => '0');
    variable r4751 : std_logic_vector(0 to 0) := (others => '0');
    variable r4750 : std_logic_vector(0 to 0) := (others => '0');
    variable r4749 : std_logic_vector(0 to 0) := (others => '0');
    variable r4748 : std_logic_vector(0 to 0) := (others => '0');
    variable r4747 : std_logic_vector(0 to 0) := (others => '0');
    variable r4746 : std_logic_vector(0 to 0) := (others => '0');
    variable r4745 : std_logic_vector(0 to 0) := (others => '0');
    variable r4744 : std_logic_vector(0 to 0) := (others => '0');
    variable r4743 : std_logic_vector(0 to 0) := (others => '0');
    variable r4742 : std_logic_vector(0 to 0) := (others => '0');
    variable r4741 : std_logic_vector(0 to 0) := (others => '0');
    variable r4740 : std_logic_vector(0 to 0) := (others => '0');
    variable r4739 : std_logic_vector(0 to 0) := (others => '0');
    variable r4738 : std_logic_vector(0 to 0) := (others => '0');
    variable r4737 : std_logic_vector(0 to 0) := (others => '0');
    variable r4736 : std_logic_vector(0 to 0) := (others => '0');
    variable r4735 : std_logic_vector(0 to 0) := (others => '0');
    variable r4734 : std_logic_vector(0 to 0) := (others => '0');
    variable r4733 : std_logic_vector(0 to 0) := (others => '0');
    variable r4732 : std_logic_vector(0 to 0) := (others => '0');
    variable r4731 : std_logic_vector(0 to 0) := (others => '0');
    variable r4730 : std_logic_vector(0 to 0) := (others => '0');
    variable r4729 : std_logic_vector(0 to 0) := (others => '0');
    variable r4728 : std_logic_vector(0 to 0) := (others => '0');
    variable r4727 : std_logic_vector(0 to 0) := (others => '0');
    variable r4726 : std_logic_vector(0 to 0) := (others => '0');
    variable r4725 : std_logic_vector(0 to 0) := (others => '0');
    variable r4724 : std_logic_vector(0 to 0) := (others => '0');
    variable r4723 : std_logic_vector(0 to 0) := (others => '0');
    variable r4722 : std_logic_vector(0 to 0) := (others => '0');
    variable r4721 : std_logic_vector(0 to 0) := (others => '0');
    variable r4720 : std_logic_vector(0 to 0) := (others => '0');
    variable r4719 : std_logic_vector(0 to 0) := (others => '0');
    variable r4718 : std_logic_vector(0 to 0) := (others => '0');
    variable r4717 : std_logic_vector(0 to 0) := (others => '0');
    variable r4716 : std_logic_vector(0 to 0) := (others => '0');
    variable r4715 : std_logic_vector(0 to 0) := (others => '0');
    variable r4714 : std_logic_vector(0 to 0) := (others => '0');
    variable r4713 : std_logic_vector(0 to 0) := (others => '0');
    variable r4712 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r4713 := "1";
    null;
    r4714 := (r4713);
    r4715 := "1";
    null;
    r4716 := (r4715);
    r4717 := "0";
    null;
    r4718 := (r4717);
    r4719 := "1";
    null;
    r4720 := (r4719);
    r4721 := "0";
    null;
    r4722 := (r4721);
    r4723 := "0";
    null;
    r4724 := (r4723);
    r4725 := "0";
    null;
    r4726 := (r4725);
    r4727 := "1";
    null;
    r4728 := (r4727);
    r4729 := "1";
    null;
    r4730 := (r4729);
    r4731 := "0";
    null;
    r4732 := (r4731);
    r4733 := "0";
    null;
    r4734 := (r4733);
    r4735 := "1";
    null;
    r4736 := (r4735);
    r4737 := "0";
    null;
    r4738 := (r4737);
    r4739 := "0";
    null;
    r4740 := (r4739);
    r4741 := "1";
    null;
    r4742 := (r4741);
    r4743 := "0";
    null;
    r4744 := (r4743);
    r4745 := "1";
    null;
    r4746 := (r4745);
    r4747 := "1";
    null;
    r4748 := (r4747);
    r4749 := "1";
    null;
    r4750 := (r4749);
    r4751 := "0";
    null;
    r4752 := (r4751);
    r4753 := "1";
    null;
    r4754 := (r4753);
    r4755 := "0";
    null;
    r4756 := (r4755);
    r4757 := "0";
    null;
    r4758 := (r4757);
    r4759 := "0";
    null;
    r4760 := (r4759);
    r4761 := "0";
    null;
    r4762 := (r4761);
    r4763 := "0";
    null;
    r4764 := (r4763);
    r4765 := "0";
    null;
    r4766 := (r4765);
    r4767 := "1";
    null;
    r4768 := (r4767);
    r4769 := "1";
    null;
    r4770 := (r4769);
    r4771 := "0";
    null;
    r4772 := (r4771);
    r4773 := "0";
    null;
    r4774 := (r4773);
    r4775 := "1";
    null;
    r4776 := (r4775);
    r4712 := (r4714 & r4716 & r4718 & r4720 & r4722 & r4724 & r4726 & r4728 & r4730 & r4732 & r4734 & r4736 & r4738 & r4740 & r4742 & r4744 & r4746 & r4748 & r4750 & r4752 & r4754 & r4756 & r4758 & r4760 & r4762 & r4764 & r4766 & r4768 & r4770 & r4772 & r4774 & r4776);
    return r4712;
  end rewire_MetaprogrammingRW.wd192e819_4711;
  function rewire_MetaprogrammingRW.wc76c51a3_4642 return std_logic_vector
  is
    variable r4707 : std_logic_vector(0 to 0) := (others => '0');
    variable r4706 : std_logic_vector(0 to 0) := (others => '0');
    variable r4705 : std_logic_vector(0 to 0) := (others => '0');
    variable r4704 : std_logic_vector(0 to 0) := (others => '0');
    variable r4703 : std_logic_vector(0 to 0) := (others => '0');
    variable r4702 : std_logic_vector(0 to 0) := (others => '0');
    variable r4701 : std_logic_vector(0 to 0) := (others => '0');
    variable r4700 : std_logic_vector(0 to 0) := (others => '0');
    variable r4699 : std_logic_vector(0 to 0) := (others => '0');
    variable r4698 : std_logic_vector(0 to 0) := (others => '0');
    variable r4697 : std_logic_vector(0 to 0) := (others => '0');
    variable r4696 : std_logic_vector(0 to 0) := (others => '0');
    variable r4695 : std_logic_vector(0 to 0) := (others => '0');
    variable r4694 : std_logic_vector(0 to 0) := (others => '0');
    variable r4693 : std_logic_vector(0 to 0) := (others => '0');
    variable r4692 : std_logic_vector(0 to 0) := (others => '0');
    variable r4691 : std_logic_vector(0 to 0) := (others => '0');
    variable r4690 : std_logic_vector(0 to 0) := (others => '0');
    variable r4689 : std_logic_vector(0 to 0) := (others => '0');
    variable r4688 : std_logic_vector(0 to 0) := (others => '0');
    variable r4687 : std_logic_vector(0 to 0) := (others => '0');
    variable r4686 : std_logic_vector(0 to 0) := (others => '0');
    variable r4685 : std_logic_vector(0 to 0) := (others => '0');
    variable r4684 : std_logic_vector(0 to 0) := (others => '0');
    variable r4683 : std_logic_vector(0 to 0) := (others => '0');
    variable r4682 : std_logic_vector(0 to 0) := (others => '0');
    variable r4681 : std_logic_vector(0 to 0) := (others => '0');
    variable r4680 : std_logic_vector(0 to 0) := (others => '0');
    variable r4679 : std_logic_vector(0 to 0) := (others => '0');
    variable r4678 : std_logic_vector(0 to 0) := (others => '0');
    variable r4677 : std_logic_vector(0 to 0) := (others => '0');
    variable r4676 : std_logic_vector(0 to 0) := (others => '0');
    variable r4675 : std_logic_vector(0 to 0) := (others => '0');
    variable r4674 : std_logic_vector(0 to 0) := (others => '0');
    variable r4673 : std_logic_vector(0 to 0) := (others => '0');
    variable r4672 : std_logic_vector(0 to 0) := (others => '0');
    variable r4671 : std_logic_vector(0 to 0) := (others => '0');
    variable r4670 : std_logic_vector(0 to 0) := (others => '0');
    variable r4669 : std_logic_vector(0 to 0) := (others => '0');
    variable r4668 : std_logic_vector(0 to 0) := (others => '0');
    variable r4667 : std_logic_vector(0 to 0) := (others => '0');
    variable r4666 : std_logic_vector(0 to 0) := (others => '0');
    variable r4665 : std_logic_vector(0 to 0) := (others => '0');
    variable r4664 : std_logic_vector(0 to 0) := (others => '0');
    variable r4663 : std_logic_vector(0 to 0) := (others => '0');
    variable r4662 : std_logic_vector(0 to 0) := (others => '0');
    variable r4661 : std_logic_vector(0 to 0) := (others => '0');
    variable r4660 : std_logic_vector(0 to 0) := (others => '0');
    variable r4659 : std_logic_vector(0 to 0) := (others => '0');
    variable r4658 : std_logic_vector(0 to 0) := (others => '0');
    variable r4657 : std_logic_vector(0 to 0) := (others => '0');
    variable r4656 : std_logic_vector(0 to 0) := (others => '0');
    variable r4655 : std_logic_vector(0 to 0) := (others => '0');
    variable r4654 : std_logic_vector(0 to 0) := (others => '0');
    variable r4653 : std_logic_vector(0 to 0) := (others => '0');
    variable r4652 : std_logic_vector(0 to 0) := (others => '0');
    variable r4651 : std_logic_vector(0 to 0) := (others => '0');
    variable r4650 : std_logic_vector(0 to 0) := (others => '0');
    variable r4649 : std_logic_vector(0 to 0) := (others => '0');
    variable r4648 : std_logic_vector(0 to 0) := (others => '0');
    variable r4647 : std_logic_vector(0 to 0) := (others => '0');
    variable r4646 : std_logic_vector(0 to 0) := (others => '0');
    variable r4645 : std_logic_vector(0 to 0) := (others => '0');
    variable r4644 : std_logic_vector(0 to 0) := (others => '0');
    variable r4643 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r4644 := "1";
    null;
    r4645 := (r4644);
    r4646 := "1";
    null;
    r4647 := (r4646);
    r4648 := "0";
    null;
    r4649 := (r4648);
    r4650 := "0";
    null;
    r4651 := (r4650);
    r4652 := "0";
    null;
    r4653 := (r4652);
    r4654 := "1";
    null;
    r4655 := (r4654);
    r4656 := "1";
    null;
    r4657 := (r4656);
    r4658 := "1";
    null;
    r4659 := (r4658);
    r4660 := "0";
    null;
    r4661 := (r4660);
    r4662 := "1";
    null;
    r4663 := (r4662);
    r4664 := "1";
    null;
    r4665 := (r4664);
    r4666 := "0";
    null;
    r4667 := (r4666);
    r4668 := "1";
    null;
    r4669 := (r4668);
    r4670 := "1";
    null;
    r4671 := (r4670);
    r4672 := "0";
    null;
    r4673 := (r4672);
    r4674 := "0";
    null;
    r4675 := (r4674);
    r4676 := "0";
    null;
    r4677 := (r4676);
    r4678 := "1";
    null;
    r4679 := (r4678);
    r4680 := "0";
    null;
    r4681 := (r4680);
    r4682 := "1";
    null;
    r4683 := (r4682);
    r4684 := "0";
    null;
    r4685 := (r4684);
    r4686 := "0";
    null;
    r4687 := (r4686);
    r4688 := "0";
    null;
    r4689 := (r4688);
    r4690 := "1";
    null;
    r4691 := (r4690);
    r4692 := "1";
    null;
    r4693 := (r4692);
    r4694 := "0";
    null;
    r4695 := (r4694);
    r4696 := "1";
    null;
    r4697 := (r4696);
    r4698 := "0";
    null;
    r4699 := (r4698);
    r4700 := "0";
    null;
    r4701 := (r4700);
    r4702 := "0";
    null;
    r4703 := (r4702);
    r4704 := "1";
    null;
    r4705 := (r4704);
    r4706 := "1";
    null;
    r4707 := (r4706);
    r4643 := (r4645 & r4647 & r4649 & r4651 & r4653 & r4655 & r4657 & r4659 & r4661 & r4663 & r4665 & r4667 & r4669 & r4671 & r4673 & r4675 & r4677 & r4679 & r4681 & r4683 & r4685 & r4687 & r4689 & r4691 & r4693 & r4695 & r4697 & r4699 & r4701 & r4703 & r4705 & r4707);
    return r4643;
  end rewire_MetaprogrammingRW.wc76c51a3_4642;
  function rewire_MetaprogrammingRW.wc24b8b70_4573 return std_logic_vector
  is
    variable r4638 : std_logic_vector(0 to 0) := (others => '0');
    variable r4637 : std_logic_vector(0 to 0) := (others => '0');
    variable r4636 : std_logic_vector(0 to 0) := (others => '0');
    variable r4635 : std_logic_vector(0 to 0) := (others => '0');
    variable r4634 : std_logic_vector(0 to 0) := (others => '0');
    variable r4633 : std_logic_vector(0 to 0) := (others => '0');
    variable r4632 : std_logic_vector(0 to 0) := (others => '0');
    variable r4631 : std_logic_vector(0 to 0) := (others => '0');
    variable r4630 : std_logic_vector(0 to 0) := (others => '0');
    variable r4629 : std_logic_vector(0 to 0) := (others => '0');
    variable r4628 : std_logic_vector(0 to 0) := (others => '0');
    variable r4627 : std_logic_vector(0 to 0) := (others => '0');
    variable r4626 : std_logic_vector(0 to 0) := (others => '0');
    variable r4625 : std_logic_vector(0 to 0) := (others => '0');
    variable r4624 : std_logic_vector(0 to 0) := (others => '0');
    variable r4623 : std_logic_vector(0 to 0) := (others => '0');
    variable r4622 : std_logic_vector(0 to 0) := (others => '0');
    variable r4621 : std_logic_vector(0 to 0) := (others => '0');
    variable r4620 : std_logic_vector(0 to 0) := (others => '0');
    variable r4619 : std_logic_vector(0 to 0) := (others => '0');
    variable r4618 : std_logic_vector(0 to 0) := (others => '0');
    variable r4617 : std_logic_vector(0 to 0) := (others => '0');
    variable r4616 : std_logic_vector(0 to 0) := (others => '0');
    variable r4615 : std_logic_vector(0 to 0) := (others => '0');
    variable r4614 : std_logic_vector(0 to 0) := (others => '0');
    variable r4613 : std_logic_vector(0 to 0) := (others => '0');
    variable r4612 : std_logic_vector(0 to 0) := (others => '0');
    variable r4611 : std_logic_vector(0 to 0) := (others => '0');
    variable r4610 : std_logic_vector(0 to 0) := (others => '0');
    variable r4609 : std_logic_vector(0 to 0) := (others => '0');
    variable r4608 : std_logic_vector(0 to 0) := (others => '0');
    variable r4607 : std_logic_vector(0 to 0) := (others => '0');
    variable r4606 : std_logic_vector(0 to 0) := (others => '0');
    variable r4605 : std_logic_vector(0 to 0) := (others => '0');
    variable r4604 : std_logic_vector(0 to 0) := (others => '0');
    variable r4603 : std_logic_vector(0 to 0) := (others => '0');
    variable r4602 : std_logic_vector(0 to 0) := (others => '0');
    variable r4601 : std_logic_vector(0 to 0) := (others => '0');
    variable r4600 : std_logic_vector(0 to 0) := (others => '0');
    variable r4599 : std_logic_vector(0 to 0) := (others => '0');
    variable r4598 : std_logic_vector(0 to 0) := (others => '0');
    variable r4597 : std_logic_vector(0 to 0) := (others => '0');
    variable r4596 : std_logic_vector(0 to 0) := (others => '0');
    variable r4595 : std_logic_vector(0 to 0) := (others => '0');
    variable r4594 : std_logic_vector(0 to 0) := (others => '0');
    variable r4593 : std_logic_vector(0 to 0) := (others => '0');
    variable r4592 : std_logic_vector(0 to 0) := (others => '0');
    variable r4591 : std_logic_vector(0 to 0) := (others => '0');
    variable r4590 : std_logic_vector(0 to 0) := (others => '0');
    variable r4589 : std_logic_vector(0 to 0) := (others => '0');
    variable r4588 : std_logic_vector(0 to 0) := (others => '0');
    variable r4587 : std_logic_vector(0 to 0) := (others => '0');
    variable r4586 : std_logic_vector(0 to 0) := (others => '0');
    variable r4585 : std_logic_vector(0 to 0) := (others => '0');
    variable r4584 : std_logic_vector(0 to 0) := (others => '0');
    variable r4583 : std_logic_vector(0 to 0) := (others => '0');
    variable r4582 : std_logic_vector(0 to 0) := (others => '0');
    variable r4581 : std_logic_vector(0 to 0) := (others => '0');
    variable r4580 : std_logic_vector(0 to 0) := (others => '0');
    variable r4579 : std_logic_vector(0 to 0) := (others => '0');
    variable r4578 : std_logic_vector(0 to 0) := (others => '0');
    variable r4577 : std_logic_vector(0 to 0) := (others => '0');
    variable r4576 : std_logic_vector(0 to 0) := (others => '0');
    variable r4575 : std_logic_vector(0 to 0) := (others => '0');
    variable r4574 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r4575 := "1";
    null;
    r4576 := (r4575);
    r4577 := "1";
    null;
    r4578 := (r4577);
    r4579 := "0";
    null;
    r4580 := (r4579);
    r4581 := "0";
    null;
    r4582 := (r4581);
    r4583 := "0";
    null;
    r4584 := (r4583);
    r4585 := "0";
    null;
    r4586 := (r4585);
    r4587 := "1";
    null;
    r4588 := (r4587);
    r4589 := "0";
    null;
    r4590 := (r4589);
    r4591 := "0";
    null;
    r4592 := (r4591);
    r4593 := "1";
    null;
    r4594 := (r4593);
    r4595 := "0";
    null;
    r4596 := (r4595);
    r4597 := "0";
    null;
    r4598 := (r4597);
    r4599 := "1";
    null;
    r4600 := (r4599);
    r4601 := "0";
    null;
    r4602 := (r4601);
    r4603 := "1";
    null;
    r4604 := (r4603);
    r4605 := "1";
    null;
    r4606 := (r4605);
    r4607 := "1";
    null;
    r4608 := (r4607);
    r4609 := "0";
    null;
    r4610 := (r4609);
    r4611 := "0";
    null;
    r4612 := (r4611);
    r4613 := "0";
    null;
    r4614 := (r4613);
    r4615 := "1";
    null;
    r4616 := (r4615);
    r4617 := "0";
    null;
    r4618 := (r4617);
    r4619 := "1";
    null;
    r4620 := (r4619);
    r4621 := "1";
    null;
    r4622 := (r4621);
    r4623 := "0";
    null;
    r4624 := (r4623);
    r4625 := "1";
    null;
    r4626 := (r4625);
    r4627 := "1";
    null;
    r4628 := (r4627);
    r4629 := "1";
    null;
    r4630 := (r4629);
    r4631 := "0";
    null;
    r4632 := (r4631);
    r4633 := "0";
    null;
    r4634 := (r4633);
    r4635 := "0";
    null;
    r4636 := (r4635);
    r4637 := "0";
    null;
    r4638 := (r4637);
    r4574 := (r4576 & r4578 & r4580 & r4582 & r4584 & r4586 & r4588 & r4590 & r4592 & r4594 & r4596 & r4598 & r4600 & r4602 & r4604 & r4606 & r4608 & r4610 & r4612 & r4614 & r4616 & r4618 & r4620 & r4622 & r4624 & r4626 & r4628 & r4630 & r4632 & r4634 & r4636 & r4638);
    return r4574;
  end rewire_MetaprogrammingRW.wc24b8b70_4573;
  function rewire_MetaprogrammingRW.wa81a664b_4504 return std_logic_vector
  is
    variable r4569 : std_logic_vector(0 to 0) := (others => '0');
    variable r4568 : std_logic_vector(0 to 0) := (others => '0');
    variable r4567 : std_logic_vector(0 to 0) := (others => '0');
    variable r4566 : std_logic_vector(0 to 0) := (others => '0');
    variable r4565 : std_logic_vector(0 to 0) := (others => '0');
    variable r4564 : std_logic_vector(0 to 0) := (others => '0');
    variable r4563 : std_logic_vector(0 to 0) := (others => '0');
    variable r4562 : std_logic_vector(0 to 0) := (others => '0');
    variable r4561 : std_logic_vector(0 to 0) := (others => '0');
    variable r4560 : std_logic_vector(0 to 0) := (others => '0');
    variable r4559 : std_logic_vector(0 to 0) := (others => '0');
    variable r4558 : std_logic_vector(0 to 0) := (others => '0');
    variable r4557 : std_logic_vector(0 to 0) := (others => '0');
    variable r4556 : std_logic_vector(0 to 0) := (others => '0');
    variable r4555 : std_logic_vector(0 to 0) := (others => '0');
    variable r4554 : std_logic_vector(0 to 0) := (others => '0');
    variable r4553 : std_logic_vector(0 to 0) := (others => '0');
    variable r4552 : std_logic_vector(0 to 0) := (others => '0');
    variable r4551 : std_logic_vector(0 to 0) := (others => '0');
    variable r4550 : std_logic_vector(0 to 0) := (others => '0');
    variable r4549 : std_logic_vector(0 to 0) := (others => '0');
    variable r4548 : std_logic_vector(0 to 0) := (others => '0');
    variable r4547 : std_logic_vector(0 to 0) := (others => '0');
    variable r4546 : std_logic_vector(0 to 0) := (others => '0');
    variable r4545 : std_logic_vector(0 to 0) := (others => '0');
    variable r4544 : std_logic_vector(0 to 0) := (others => '0');
    variable r4543 : std_logic_vector(0 to 0) := (others => '0');
    variable r4542 : std_logic_vector(0 to 0) := (others => '0');
    variable r4541 : std_logic_vector(0 to 0) := (others => '0');
    variable r4540 : std_logic_vector(0 to 0) := (others => '0');
    variable r4539 : std_logic_vector(0 to 0) := (others => '0');
    variable r4538 : std_logic_vector(0 to 0) := (others => '0');
    variable r4537 : std_logic_vector(0 to 0) := (others => '0');
    variable r4536 : std_logic_vector(0 to 0) := (others => '0');
    variable r4535 : std_logic_vector(0 to 0) := (others => '0');
    variable r4534 : std_logic_vector(0 to 0) := (others => '0');
    variable r4533 : std_logic_vector(0 to 0) := (others => '0');
    variable r4532 : std_logic_vector(0 to 0) := (others => '0');
    variable r4531 : std_logic_vector(0 to 0) := (others => '0');
    variable r4530 : std_logic_vector(0 to 0) := (others => '0');
    variable r4529 : std_logic_vector(0 to 0) := (others => '0');
    variable r4528 : std_logic_vector(0 to 0) := (others => '0');
    variable r4527 : std_logic_vector(0 to 0) := (others => '0');
    variable r4526 : std_logic_vector(0 to 0) := (others => '0');
    variable r4525 : std_logic_vector(0 to 0) := (others => '0');
    variable r4524 : std_logic_vector(0 to 0) := (others => '0');
    variable r4523 : std_logic_vector(0 to 0) := (others => '0');
    variable r4522 : std_logic_vector(0 to 0) := (others => '0');
    variable r4521 : std_logic_vector(0 to 0) := (others => '0');
    variable r4520 : std_logic_vector(0 to 0) := (others => '0');
    variable r4519 : std_logic_vector(0 to 0) := (others => '0');
    variable r4518 : std_logic_vector(0 to 0) := (others => '0');
    variable r4517 : std_logic_vector(0 to 0) := (others => '0');
    variable r4516 : std_logic_vector(0 to 0) := (others => '0');
    variable r4515 : std_logic_vector(0 to 0) := (others => '0');
    variable r4514 : std_logic_vector(0 to 0) := (others => '0');
    variable r4513 : std_logic_vector(0 to 0) := (others => '0');
    variable r4512 : std_logic_vector(0 to 0) := (others => '0');
    variable r4511 : std_logic_vector(0 to 0) := (others => '0');
    variable r4510 : std_logic_vector(0 to 0) := (others => '0');
    variable r4509 : std_logic_vector(0 to 0) := (others => '0');
    variable r4508 : std_logic_vector(0 to 0) := (others => '0');
    variable r4507 : std_logic_vector(0 to 0) := (others => '0');
    variable r4506 : std_logic_vector(0 to 0) := (others => '0');
    variable r4505 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r4506 := "1";
    null;
    r4507 := (r4506);
    r4508 := "0";
    null;
    r4509 := (r4508);
    r4510 := "1";
    null;
    r4511 := (r4510);
    r4512 := "0";
    null;
    r4513 := (r4512);
    r4514 := "1";
    null;
    r4515 := (r4514);
    r4516 := "0";
    null;
    r4517 := (r4516);
    r4518 := "0";
    null;
    r4519 := (r4518);
    r4520 := "0";
    null;
    r4521 := (r4520);
    r4522 := "0";
    null;
    r4523 := (r4522);
    r4524 := "0";
    null;
    r4525 := (r4524);
    r4526 := "0";
    null;
    r4527 := (r4526);
    r4528 := "1";
    null;
    r4529 := (r4528);
    r4530 := "1";
    null;
    r4531 := (r4530);
    r4532 := "0";
    null;
    r4533 := (r4532);
    r4534 := "1";
    null;
    r4535 := (r4534);
    r4536 := "0";
    null;
    r4537 := (r4536);
    r4538 := "0";
    null;
    r4539 := (r4538);
    r4540 := "1";
    null;
    r4541 := (r4540);
    r4542 := "1";
    null;
    r4543 := (r4542);
    r4544 := "0";
    null;
    r4545 := (r4544);
    r4546 := "0";
    null;
    r4547 := (r4546);
    r4548 := "1";
    null;
    r4549 := (r4548);
    r4550 := "1";
    null;
    r4551 := (r4550);
    r4552 := "0";
    null;
    r4553 := (r4552);
    r4554 := "0";
    null;
    r4555 := (r4554);
    r4556 := "1";
    null;
    r4557 := (r4556);
    r4558 := "0";
    null;
    r4559 := (r4558);
    r4560 := "0";
    null;
    r4561 := (r4560);
    r4562 := "1";
    null;
    r4563 := (r4562);
    r4564 := "0";
    null;
    r4565 := (r4564);
    r4566 := "1";
    null;
    r4567 := (r4566);
    r4568 := "1";
    null;
    r4569 := (r4568);
    r4505 := (r4507 & r4509 & r4511 & r4513 & r4515 & r4517 & r4519 & r4521 & r4523 & r4525 & r4527 & r4529 & r4531 & r4533 & r4535 & r4537 & r4539 & r4541 & r4543 & r4545 & r4547 & r4549 & r4551 & r4553 & r4555 & r4557 & r4559 & r4561 & r4563 & r4565 & r4567 & r4569);
    return r4505;
  end rewire_MetaprogrammingRW.wa81a664b_4504;
  function rewire_MetaprogrammingRW.wa2bfe8a1_4435 return std_logic_vector
  is
    variable r4500 : std_logic_vector(0 to 0) := (others => '0');
    variable r4499 : std_logic_vector(0 to 0) := (others => '0');
    variable r4498 : std_logic_vector(0 to 0) := (others => '0');
    variable r4497 : std_logic_vector(0 to 0) := (others => '0');
    variable r4496 : std_logic_vector(0 to 0) := (others => '0');
    variable r4495 : std_logic_vector(0 to 0) := (others => '0');
    variable r4494 : std_logic_vector(0 to 0) := (others => '0');
    variable r4493 : std_logic_vector(0 to 0) := (others => '0');
    variable r4492 : std_logic_vector(0 to 0) := (others => '0');
    variable r4491 : std_logic_vector(0 to 0) := (others => '0');
    variable r4490 : std_logic_vector(0 to 0) := (others => '0');
    variable r4489 : std_logic_vector(0 to 0) := (others => '0');
    variable r4488 : std_logic_vector(0 to 0) := (others => '0');
    variable r4487 : std_logic_vector(0 to 0) := (others => '0');
    variable r4486 : std_logic_vector(0 to 0) := (others => '0');
    variable r4485 : std_logic_vector(0 to 0) := (others => '0');
    variable r4484 : std_logic_vector(0 to 0) := (others => '0');
    variable r4483 : std_logic_vector(0 to 0) := (others => '0');
    variable r4482 : std_logic_vector(0 to 0) := (others => '0');
    variable r4481 : std_logic_vector(0 to 0) := (others => '0');
    variable r4480 : std_logic_vector(0 to 0) := (others => '0');
    variable r4479 : std_logic_vector(0 to 0) := (others => '0');
    variable r4478 : std_logic_vector(0 to 0) := (others => '0');
    variable r4477 : std_logic_vector(0 to 0) := (others => '0');
    variable r4476 : std_logic_vector(0 to 0) := (others => '0');
    variable r4475 : std_logic_vector(0 to 0) := (others => '0');
    variable r4474 : std_logic_vector(0 to 0) := (others => '0');
    variable r4473 : std_logic_vector(0 to 0) := (others => '0');
    variable r4472 : std_logic_vector(0 to 0) := (others => '0');
    variable r4471 : std_logic_vector(0 to 0) := (others => '0');
    variable r4470 : std_logic_vector(0 to 0) := (others => '0');
    variable r4469 : std_logic_vector(0 to 0) := (others => '0');
    variable r4468 : std_logic_vector(0 to 0) := (others => '0');
    variable r4467 : std_logic_vector(0 to 0) := (others => '0');
    variable r4466 : std_logic_vector(0 to 0) := (others => '0');
    variable r4465 : std_logic_vector(0 to 0) := (others => '0');
    variable r4464 : std_logic_vector(0 to 0) := (others => '0');
    variable r4463 : std_logic_vector(0 to 0) := (others => '0');
    variable r4462 : std_logic_vector(0 to 0) := (others => '0');
    variable r4461 : std_logic_vector(0 to 0) := (others => '0');
    variable r4460 : std_logic_vector(0 to 0) := (others => '0');
    variable r4459 : std_logic_vector(0 to 0) := (others => '0');
    variable r4458 : std_logic_vector(0 to 0) := (others => '0');
    variable r4457 : std_logic_vector(0 to 0) := (others => '0');
    variable r4456 : std_logic_vector(0 to 0) := (others => '0');
    variable r4455 : std_logic_vector(0 to 0) := (others => '0');
    variable r4454 : std_logic_vector(0 to 0) := (others => '0');
    variable r4453 : std_logic_vector(0 to 0) := (others => '0');
    variable r4452 : std_logic_vector(0 to 0) := (others => '0');
    variable r4451 : std_logic_vector(0 to 0) := (others => '0');
    variable r4450 : std_logic_vector(0 to 0) := (others => '0');
    variable r4449 : std_logic_vector(0 to 0) := (others => '0');
    variable r4448 : std_logic_vector(0 to 0) := (others => '0');
    variable r4447 : std_logic_vector(0 to 0) := (others => '0');
    variable r4446 : std_logic_vector(0 to 0) := (others => '0');
    variable r4445 : std_logic_vector(0 to 0) := (others => '0');
    variable r4444 : std_logic_vector(0 to 0) := (others => '0');
    variable r4443 : std_logic_vector(0 to 0) := (others => '0');
    variable r4442 : std_logic_vector(0 to 0) := (others => '0');
    variable r4441 : std_logic_vector(0 to 0) := (others => '0');
    variable r4440 : std_logic_vector(0 to 0) := (others => '0');
    variable r4439 : std_logic_vector(0 to 0) := (others => '0');
    variable r4438 : std_logic_vector(0 to 0) := (others => '0');
    variable r4437 : std_logic_vector(0 to 0) := (others => '0');
    variable r4436 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r4437 := "1";
    null;
    r4438 := (r4437);
    r4439 := "0";
    null;
    r4440 := (r4439);
    r4441 := "1";
    null;
    r4442 := (r4441);
    r4443 := "0";
    null;
    r4444 := (r4443);
    r4445 := "0";
    null;
    r4446 := (r4445);
    r4447 := "0";
    null;
    r4448 := (r4447);
    r4449 := "1";
    null;
    r4450 := (r4449);
    r4451 := "0";
    null;
    r4452 := (r4451);
    r4453 := "1";
    null;
    r4454 := (r4453);
    r4455 := "0";
    null;
    r4456 := (r4455);
    r4457 := "1";
    null;
    r4458 := (r4457);
    r4459 := "1";
    null;
    r4460 := (r4459);
    r4461 := "1";
    null;
    r4462 := (r4461);
    r4463 := "1";
    null;
    r4464 := (r4463);
    r4465 := "1";
    null;
    r4466 := (r4465);
    r4467 := "1";
    null;
    r4468 := (r4467);
    r4469 := "1";
    null;
    r4470 := (r4469);
    r4471 := "1";
    null;
    r4472 := (r4471);
    r4473 := "1";
    null;
    r4474 := (r4473);
    r4475 := "0";
    null;
    r4476 := (r4475);
    r4477 := "1";
    null;
    r4478 := (r4477);
    r4479 := "0";
    null;
    r4480 := (r4479);
    r4481 := "0";
    null;
    r4482 := (r4481);
    r4483 := "0";
    null;
    r4484 := (r4483);
    r4485 := "1";
    null;
    r4486 := (r4485);
    r4487 := "0";
    null;
    r4488 := (r4487);
    r4489 := "1";
    null;
    r4490 := (r4489);
    r4491 := "0";
    null;
    r4492 := (r4491);
    r4493 := "0";
    null;
    r4494 := (r4493);
    r4495 := "0";
    null;
    r4496 := (r4495);
    r4497 := "0";
    null;
    r4498 := (r4497);
    r4499 := "1";
    null;
    r4500 := (r4499);
    r4436 := (r4438 & r4440 & r4442 & r4444 & r4446 & r4448 & r4450 & r4452 & r4454 & r4456 & r4458 & r4460 & r4462 & r4464 & r4466 & r4468 & r4470 & r4472 & r4474 & r4476 & r4478 & r4480 & r4482 & r4484 & r4486 & r4488 & r4490 & r4492 & r4494 & r4496 & r4498 & r4500);
    return r4436;
  end rewire_MetaprogrammingRW.wa2bfe8a1_4435;
  function rewire_MetaprogrammingRW.w92722c85_4366 return std_logic_vector
  is
    variable r4431 : std_logic_vector(0 to 0) := (others => '0');
    variable r4430 : std_logic_vector(0 to 0) := (others => '0');
    variable r4429 : std_logic_vector(0 to 0) := (others => '0');
    variable r4428 : std_logic_vector(0 to 0) := (others => '0');
    variable r4427 : std_logic_vector(0 to 0) := (others => '0');
    variable r4426 : std_logic_vector(0 to 0) := (others => '0');
    variable r4425 : std_logic_vector(0 to 0) := (others => '0');
    variable r4424 : std_logic_vector(0 to 0) := (others => '0');
    variable r4423 : std_logic_vector(0 to 0) := (others => '0');
    variable r4422 : std_logic_vector(0 to 0) := (others => '0');
    variable r4421 : std_logic_vector(0 to 0) := (others => '0');
    variable r4420 : std_logic_vector(0 to 0) := (others => '0');
    variable r4419 : std_logic_vector(0 to 0) := (others => '0');
    variable r4418 : std_logic_vector(0 to 0) := (others => '0');
    variable r4417 : std_logic_vector(0 to 0) := (others => '0');
    variable r4416 : std_logic_vector(0 to 0) := (others => '0');
    variable r4415 : std_logic_vector(0 to 0) := (others => '0');
    variable r4414 : std_logic_vector(0 to 0) := (others => '0');
    variable r4413 : std_logic_vector(0 to 0) := (others => '0');
    variable r4412 : std_logic_vector(0 to 0) := (others => '0');
    variable r4411 : std_logic_vector(0 to 0) := (others => '0');
    variable r4410 : std_logic_vector(0 to 0) := (others => '0');
    variable r4409 : std_logic_vector(0 to 0) := (others => '0');
    variable r4408 : std_logic_vector(0 to 0) := (others => '0');
    variable r4407 : std_logic_vector(0 to 0) := (others => '0');
    variable r4406 : std_logic_vector(0 to 0) := (others => '0');
    variable r4405 : std_logic_vector(0 to 0) := (others => '0');
    variable r4404 : std_logic_vector(0 to 0) := (others => '0');
    variable r4403 : std_logic_vector(0 to 0) := (others => '0');
    variable r4402 : std_logic_vector(0 to 0) := (others => '0');
    variable r4401 : std_logic_vector(0 to 0) := (others => '0');
    variable r4400 : std_logic_vector(0 to 0) := (others => '0');
    variable r4399 : std_logic_vector(0 to 0) := (others => '0');
    variable r4398 : std_logic_vector(0 to 0) := (others => '0');
    variable r4397 : std_logic_vector(0 to 0) := (others => '0');
    variable r4396 : std_logic_vector(0 to 0) := (others => '0');
    variable r4395 : std_logic_vector(0 to 0) := (others => '0');
    variable r4394 : std_logic_vector(0 to 0) := (others => '0');
    variable r4393 : std_logic_vector(0 to 0) := (others => '0');
    variable r4392 : std_logic_vector(0 to 0) := (others => '0');
    variable r4391 : std_logic_vector(0 to 0) := (others => '0');
    variable r4390 : std_logic_vector(0 to 0) := (others => '0');
    variable r4389 : std_logic_vector(0 to 0) := (others => '0');
    variable r4388 : std_logic_vector(0 to 0) := (others => '0');
    variable r4387 : std_logic_vector(0 to 0) := (others => '0');
    variable r4386 : std_logic_vector(0 to 0) := (others => '0');
    variable r4385 : std_logic_vector(0 to 0) := (others => '0');
    variable r4384 : std_logic_vector(0 to 0) := (others => '0');
    variable r4383 : std_logic_vector(0 to 0) := (others => '0');
    variable r4382 : std_logic_vector(0 to 0) := (others => '0');
    variable r4381 : std_logic_vector(0 to 0) := (others => '0');
    variable r4380 : std_logic_vector(0 to 0) := (others => '0');
    variable r4379 : std_logic_vector(0 to 0) := (others => '0');
    variable r4378 : std_logic_vector(0 to 0) := (others => '0');
    variable r4377 : std_logic_vector(0 to 0) := (others => '0');
    variable r4376 : std_logic_vector(0 to 0) := (others => '0');
    variable r4375 : std_logic_vector(0 to 0) := (others => '0');
    variable r4374 : std_logic_vector(0 to 0) := (others => '0');
    variable r4373 : std_logic_vector(0 to 0) := (others => '0');
    variable r4372 : std_logic_vector(0 to 0) := (others => '0');
    variable r4371 : std_logic_vector(0 to 0) := (others => '0');
    variable r4370 : std_logic_vector(0 to 0) := (others => '0');
    variable r4369 : std_logic_vector(0 to 0) := (others => '0');
    variable r4368 : std_logic_vector(0 to 0) := (others => '0');
    variable r4367 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r4368 := "1";
    null;
    r4369 := (r4368);
    r4370 := "0";
    null;
    r4371 := (r4370);
    r4372 := "0";
    null;
    r4373 := (r4372);
    r4374 := "1";
    null;
    r4375 := (r4374);
    r4376 := "0";
    null;
    r4377 := (r4376);
    r4378 := "0";
    null;
    r4379 := (r4378);
    r4380 := "1";
    null;
    r4381 := (r4380);
    r4382 := "0";
    null;
    r4383 := (r4382);
    r4384 := "0";
    null;
    r4385 := (r4384);
    r4386 := "1";
    null;
    r4387 := (r4386);
    r4388 := "1";
    null;
    r4389 := (r4388);
    r4390 := "1";
    null;
    r4391 := (r4390);
    r4392 := "0";
    null;
    r4393 := (r4392);
    r4394 := "0";
    null;
    r4395 := (r4394);
    r4396 := "1";
    null;
    r4397 := (r4396);
    r4398 := "0";
    null;
    r4399 := (r4398);
    r4400 := "0";
    null;
    r4401 := (r4400);
    r4402 := "0";
    null;
    r4403 := (r4402);
    r4404 := "1";
    null;
    r4405 := (r4404);
    r4406 := "0";
    null;
    r4407 := (r4406);
    r4408 := "1";
    null;
    r4409 := (r4408);
    r4410 := "1";
    null;
    r4411 := (r4410);
    r4412 := "0";
    null;
    r4413 := (r4412);
    r4414 := "0";
    null;
    r4415 := (r4414);
    r4416 := "1";
    null;
    r4417 := (r4416);
    r4418 := "0";
    null;
    r4419 := (r4418);
    r4420 := "0";
    null;
    r4421 := (r4420);
    r4422 := "0";
    null;
    r4423 := (r4422);
    r4424 := "0";
    null;
    r4425 := (r4424);
    r4426 := "1";
    null;
    r4427 := (r4426);
    r4428 := "0";
    null;
    r4429 := (r4428);
    r4430 := "1";
    null;
    r4431 := (r4430);
    r4367 := (r4369 & r4371 & r4373 & r4375 & r4377 & r4379 & r4381 & r4383 & r4385 & r4387 & r4389 & r4391 & r4393 & r4395 & r4397 & r4399 & r4401 & r4403 & r4405 & r4407 & r4409 & r4411 & r4413 & r4415 & r4417 & r4419 & r4421 & r4423 & r4425 & r4427 & r4429 & r4431);
    return r4367;
  end rewire_MetaprogrammingRW.w92722c85_4366;
  function rewire_MetaprogrammingRW.w81c2c92e_4297 return std_logic_vector
  is
    variable r4362 : std_logic_vector(0 to 0) := (others => '0');
    variable r4361 : std_logic_vector(0 to 0) := (others => '0');
    variable r4360 : std_logic_vector(0 to 0) := (others => '0');
    variable r4359 : std_logic_vector(0 to 0) := (others => '0');
    variable r4358 : std_logic_vector(0 to 0) := (others => '0');
    variable r4357 : std_logic_vector(0 to 0) := (others => '0');
    variable r4356 : std_logic_vector(0 to 0) := (others => '0');
    variable r4355 : std_logic_vector(0 to 0) := (others => '0');
    variable r4354 : std_logic_vector(0 to 0) := (others => '0');
    variable r4353 : std_logic_vector(0 to 0) := (others => '0');
    variable r4352 : std_logic_vector(0 to 0) := (others => '0');
    variable r4351 : std_logic_vector(0 to 0) := (others => '0');
    variable r4350 : std_logic_vector(0 to 0) := (others => '0');
    variable r4349 : std_logic_vector(0 to 0) := (others => '0');
    variable r4348 : std_logic_vector(0 to 0) := (others => '0');
    variable r4347 : std_logic_vector(0 to 0) := (others => '0');
    variable r4346 : std_logic_vector(0 to 0) := (others => '0');
    variable r4345 : std_logic_vector(0 to 0) := (others => '0');
    variable r4344 : std_logic_vector(0 to 0) := (others => '0');
    variable r4343 : std_logic_vector(0 to 0) := (others => '0');
    variable r4342 : std_logic_vector(0 to 0) := (others => '0');
    variable r4341 : std_logic_vector(0 to 0) := (others => '0');
    variable r4340 : std_logic_vector(0 to 0) := (others => '0');
    variable r4339 : std_logic_vector(0 to 0) := (others => '0');
    variable r4338 : std_logic_vector(0 to 0) := (others => '0');
    variable r4337 : std_logic_vector(0 to 0) := (others => '0');
    variable r4336 : std_logic_vector(0 to 0) := (others => '0');
    variable r4335 : std_logic_vector(0 to 0) := (others => '0');
    variable r4334 : std_logic_vector(0 to 0) := (others => '0');
    variable r4333 : std_logic_vector(0 to 0) := (others => '0');
    variable r4332 : std_logic_vector(0 to 0) := (others => '0');
    variable r4331 : std_logic_vector(0 to 0) := (others => '0');
    variable r4330 : std_logic_vector(0 to 0) := (others => '0');
    variable r4329 : std_logic_vector(0 to 0) := (others => '0');
    variable r4328 : std_logic_vector(0 to 0) := (others => '0');
    variable r4327 : std_logic_vector(0 to 0) := (others => '0');
    variable r4326 : std_logic_vector(0 to 0) := (others => '0');
    variable r4325 : std_logic_vector(0 to 0) := (others => '0');
    variable r4324 : std_logic_vector(0 to 0) := (others => '0');
    variable r4323 : std_logic_vector(0 to 0) := (others => '0');
    variable r4322 : std_logic_vector(0 to 0) := (others => '0');
    variable r4321 : std_logic_vector(0 to 0) := (others => '0');
    variable r4320 : std_logic_vector(0 to 0) := (others => '0');
    variable r4319 : std_logic_vector(0 to 0) := (others => '0');
    variable r4318 : std_logic_vector(0 to 0) := (others => '0');
    variable r4317 : std_logic_vector(0 to 0) := (others => '0');
    variable r4316 : std_logic_vector(0 to 0) := (others => '0');
    variable r4315 : std_logic_vector(0 to 0) := (others => '0');
    variable r4314 : std_logic_vector(0 to 0) := (others => '0');
    variable r4313 : std_logic_vector(0 to 0) := (others => '0');
    variable r4312 : std_logic_vector(0 to 0) := (others => '0');
    variable r4311 : std_logic_vector(0 to 0) := (others => '0');
    variable r4310 : std_logic_vector(0 to 0) := (others => '0');
    variable r4309 : std_logic_vector(0 to 0) := (others => '0');
    variable r4308 : std_logic_vector(0 to 0) := (others => '0');
    variable r4307 : std_logic_vector(0 to 0) := (others => '0');
    variable r4306 : std_logic_vector(0 to 0) := (others => '0');
    variable r4305 : std_logic_vector(0 to 0) := (others => '0');
    variable r4304 : std_logic_vector(0 to 0) := (others => '0');
    variable r4303 : std_logic_vector(0 to 0) := (others => '0');
    variable r4302 : std_logic_vector(0 to 0) := (others => '0');
    variable r4301 : std_logic_vector(0 to 0) := (others => '0');
    variable r4300 : std_logic_vector(0 to 0) := (others => '0');
    variable r4299 : std_logic_vector(0 to 0) := (others => '0');
    variable r4298 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r4299 := "1";
    null;
    r4300 := (r4299);
    r4301 := "0";
    null;
    r4302 := (r4301);
    r4303 := "0";
    null;
    r4304 := (r4303);
    r4305 := "0";
    null;
    r4306 := (r4305);
    r4307 := "0";
    null;
    r4308 := (r4307);
    r4309 := "0";
    null;
    r4310 := (r4309);
    r4311 := "0";
    null;
    r4312 := (r4311);
    r4313 := "1";
    null;
    r4314 := (r4313);
    r4315 := "1";
    null;
    r4316 := (r4315);
    r4317 := "1";
    null;
    r4318 := (r4317);
    r4319 := "0";
    null;
    r4320 := (r4319);
    r4321 := "0";
    null;
    r4322 := (r4321);
    r4323 := "0";
    null;
    r4324 := (r4323);
    r4325 := "0";
    null;
    r4326 := (r4325);
    r4327 := "1";
    null;
    r4328 := (r4327);
    r4329 := "0";
    null;
    r4330 := (r4329);
    r4331 := "1";
    null;
    r4332 := (r4331);
    r4333 := "1";
    null;
    r4334 := (r4333);
    r4335 := "0";
    null;
    r4336 := (r4335);
    r4337 := "0";
    null;
    r4338 := (r4337);
    r4339 := "1";
    null;
    r4340 := (r4339);
    r4341 := "0";
    null;
    r4342 := (r4341);
    r4343 := "0";
    null;
    r4344 := (r4343);
    r4345 := "1";
    null;
    r4346 := (r4345);
    r4347 := "0";
    null;
    r4348 := (r4347);
    r4349 := "0";
    null;
    r4350 := (r4349);
    r4351 := "1";
    null;
    r4352 := (r4351);
    r4353 := "0";
    null;
    r4354 := (r4353);
    r4355 := "1";
    null;
    r4356 := (r4355);
    r4357 := "1";
    null;
    r4358 := (r4357);
    r4359 := "1";
    null;
    r4360 := (r4359);
    r4361 := "0";
    null;
    r4362 := (r4361);
    r4298 := (r4300 & r4302 & r4304 & r4306 & r4308 & r4310 & r4312 & r4314 & r4316 & r4318 & r4320 & r4322 & r4324 & r4326 & r4328 & r4330 & r4332 & r4334 & r4336 & r4338 & r4340 & r4342 & r4344 & r4346 & r4348 & r4350 & r4352 & r4354 & r4356 & r4358 & r4360 & r4362);
    return r4298;
  end rewire_MetaprogrammingRW.w81c2c92e_4297;
  function rewire_MetaprogrammingRW.w766a0abb_4228 return std_logic_vector
  is
    variable r4293 : std_logic_vector(0 to 0) := (others => '0');
    variable r4292 : std_logic_vector(0 to 0) := (others => '0');
    variable r4291 : std_logic_vector(0 to 0) := (others => '0');
    variable r4290 : std_logic_vector(0 to 0) := (others => '0');
    variable r4289 : std_logic_vector(0 to 0) := (others => '0');
    variable r4288 : std_logic_vector(0 to 0) := (others => '0');
    variable r4287 : std_logic_vector(0 to 0) := (others => '0');
    variable r4286 : std_logic_vector(0 to 0) := (others => '0');
    variable r4285 : std_logic_vector(0 to 0) := (others => '0');
    variable r4284 : std_logic_vector(0 to 0) := (others => '0');
    variable r4283 : std_logic_vector(0 to 0) := (others => '0');
    variable r4282 : std_logic_vector(0 to 0) := (others => '0');
    variable r4281 : std_logic_vector(0 to 0) := (others => '0');
    variable r4280 : std_logic_vector(0 to 0) := (others => '0');
    variable r4279 : std_logic_vector(0 to 0) := (others => '0');
    variable r4278 : std_logic_vector(0 to 0) := (others => '0');
    variable r4277 : std_logic_vector(0 to 0) := (others => '0');
    variable r4276 : std_logic_vector(0 to 0) := (others => '0');
    variable r4275 : std_logic_vector(0 to 0) := (others => '0');
    variable r4274 : std_logic_vector(0 to 0) := (others => '0');
    variable r4273 : std_logic_vector(0 to 0) := (others => '0');
    variable r4272 : std_logic_vector(0 to 0) := (others => '0');
    variable r4271 : std_logic_vector(0 to 0) := (others => '0');
    variable r4270 : std_logic_vector(0 to 0) := (others => '0');
    variable r4269 : std_logic_vector(0 to 0) := (others => '0');
    variable r4268 : std_logic_vector(0 to 0) := (others => '0');
    variable r4267 : std_logic_vector(0 to 0) := (others => '0');
    variable r4266 : std_logic_vector(0 to 0) := (others => '0');
    variable r4265 : std_logic_vector(0 to 0) := (others => '0');
    variable r4264 : std_logic_vector(0 to 0) := (others => '0');
    variable r4263 : std_logic_vector(0 to 0) := (others => '0');
    variable r4262 : std_logic_vector(0 to 0) := (others => '0');
    variable r4261 : std_logic_vector(0 to 0) := (others => '0');
    variable r4260 : std_logic_vector(0 to 0) := (others => '0');
    variable r4259 : std_logic_vector(0 to 0) := (others => '0');
    variable r4258 : std_logic_vector(0 to 0) := (others => '0');
    variable r4257 : std_logic_vector(0 to 0) := (others => '0');
    variable r4256 : std_logic_vector(0 to 0) := (others => '0');
    variable r4255 : std_logic_vector(0 to 0) := (others => '0');
    variable r4254 : std_logic_vector(0 to 0) := (others => '0');
    variable r4253 : std_logic_vector(0 to 0) := (others => '0');
    variable r4252 : std_logic_vector(0 to 0) := (others => '0');
    variable r4251 : std_logic_vector(0 to 0) := (others => '0');
    variable r4250 : std_logic_vector(0 to 0) := (others => '0');
    variable r4249 : std_logic_vector(0 to 0) := (others => '0');
    variable r4248 : std_logic_vector(0 to 0) := (others => '0');
    variable r4247 : std_logic_vector(0 to 0) := (others => '0');
    variable r4246 : std_logic_vector(0 to 0) := (others => '0');
    variable r4245 : std_logic_vector(0 to 0) := (others => '0');
    variable r4244 : std_logic_vector(0 to 0) := (others => '0');
    variable r4243 : std_logic_vector(0 to 0) := (others => '0');
    variable r4242 : std_logic_vector(0 to 0) := (others => '0');
    variable r4241 : std_logic_vector(0 to 0) := (others => '0');
    variable r4240 : std_logic_vector(0 to 0) := (others => '0');
    variable r4239 : std_logic_vector(0 to 0) := (others => '0');
    variable r4238 : std_logic_vector(0 to 0) := (others => '0');
    variable r4237 : std_logic_vector(0 to 0) := (others => '0');
    variable r4236 : std_logic_vector(0 to 0) := (others => '0');
    variable r4235 : std_logic_vector(0 to 0) := (others => '0');
    variable r4234 : std_logic_vector(0 to 0) := (others => '0');
    variable r4233 : std_logic_vector(0 to 0) := (others => '0');
    variable r4232 : std_logic_vector(0 to 0) := (others => '0');
    variable r4231 : std_logic_vector(0 to 0) := (others => '0');
    variable r4230 : std_logic_vector(0 to 0) := (others => '0');
    variable r4229 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r4230 := "0";
    null;
    r4231 := (r4230);
    r4232 := "1";
    null;
    r4233 := (r4232);
    r4234 := "1";
    null;
    r4235 := (r4234);
    r4236 := "1";
    null;
    r4237 := (r4236);
    r4238 := "0";
    null;
    r4239 := (r4238);
    r4240 := "1";
    null;
    r4241 := (r4240);
    r4242 := "1";
    null;
    r4243 := (r4242);
    r4244 := "0";
    null;
    r4245 := (r4244);
    r4246 := "0";
    null;
    r4247 := (r4246);
    r4248 := "1";
    null;
    r4249 := (r4248);
    r4250 := "1";
    null;
    r4251 := (r4250);
    r4252 := "0";
    null;
    r4253 := (r4252);
    r4254 := "1";
    null;
    r4255 := (r4254);
    r4256 := "0";
    null;
    r4257 := (r4256);
    r4258 := "1";
    null;
    r4259 := (r4258);
    r4260 := "0";
    null;
    r4261 := (r4260);
    r4262 := "0";
    null;
    r4263 := (r4262);
    r4264 := "0";
    null;
    r4265 := (r4264);
    r4266 := "0";
    null;
    r4267 := (r4266);
    r4268 := "0";
    null;
    r4269 := (r4268);
    r4270 := "1";
    null;
    r4271 := (r4270);
    r4272 := "0";
    null;
    r4273 := (r4272);
    r4274 := "1";
    null;
    r4275 := (r4274);
    r4276 := "0";
    null;
    r4277 := (r4276);
    r4278 := "1";
    null;
    r4279 := (r4278);
    r4280 := "0";
    null;
    r4281 := (r4280);
    r4282 := "1";
    null;
    r4283 := (r4282);
    r4284 := "1";
    null;
    r4285 := (r4284);
    r4286 := "1";
    null;
    r4287 := (r4286);
    r4288 := "0";
    null;
    r4289 := (r4288);
    r4290 := "1";
    null;
    r4291 := (r4290);
    r4292 := "1";
    null;
    r4293 := (r4292);
    r4229 := (r4231 & r4233 & r4235 & r4237 & r4239 & r4241 & r4243 & r4245 & r4247 & r4249 & r4251 & r4253 & r4255 & r4257 & r4259 & r4261 & r4263 & r4265 & r4267 & r4269 & r4271 & r4273 & r4275 & r4277 & r4279 & r4281 & r4283 & r4285 & r4287 & r4289 & r4291 & r4293);
    return r4229;
  end rewire_MetaprogrammingRW.w766a0abb_4228;
  function rewire_MetaprogrammingRW.w650a7354_4159 return std_logic_vector
  is
    variable r4224 : std_logic_vector(0 to 0) := (others => '0');
    variable r4223 : std_logic_vector(0 to 0) := (others => '0');
    variable r4222 : std_logic_vector(0 to 0) := (others => '0');
    variable r4221 : std_logic_vector(0 to 0) := (others => '0');
    variable r4220 : std_logic_vector(0 to 0) := (others => '0');
    variable r4219 : std_logic_vector(0 to 0) := (others => '0');
    variable r4218 : std_logic_vector(0 to 0) := (others => '0');
    variable r4217 : std_logic_vector(0 to 0) := (others => '0');
    variable r4216 : std_logic_vector(0 to 0) := (others => '0');
    variable r4215 : std_logic_vector(0 to 0) := (others => '0');
    variable r4214 : std_logic_vector(0 to 0) := (others => '0');
    variable r4213 : std_logic_vector(0 to 0) := (others => '0');
    variable r4212 : std_logic_vector(0 to 0) := (others => '0');
    variable r4211 : std_logic_vector(0 to 0) := (others => '0');
    variable r4210 : std_logic_vector(0 to 0) := (others => '0');
    variable r4209 : std_logic_vector(0 to 0) := (others => '0');
    variable r4208 : std_logic_vector(0 to 0) := (others => '0');
    variable r4207 : std_logic_vector(0 to 0) := (others => '0');
    variable r4206 : std_logic_vector(0 to 0) := (others => '0');
    variable r4205 : std_logic_vector(0 to 0) := (others => '0');
    variable r4204 : std_logic_vector(0 to 0) := (others => '0');
    variable r4203 : std_logic_vector(0 to 0) := (others => '0');
    variable r4202 : std_logic_vector(0 to 0) := (others => '0');
    variable r4201 : std_logic_vector(0 to 0) := (others => '0');
    variable r4200 : std_logic_vector(0 to 0) := (others => '0');
    variable r4199 : std_logic_vector(0 to 0) := (others => '0');
    variable r4198 : std_logic_vector(0 to 0) := (others => '0');
    variable r4197 : std_logic_vector(0 to 0) := (others => '0');
    variable r4196 : std_logic_vector(0 to 0) := (others => '0');
    variable r4195 : std_logic_vector(0 to 0) := (others => '0');
    variable r4194 : std_logic_vector(0 to 0) := (others => '0');
    variable r4193 : std_logic_vector(0 to 0) := (others => '0');
    variable r4192 : std_logic_vector(0 to 0) := (others => '0');
    variable r4191 : std_logic_vector(0 to 0) := (others => '0');
    variable r4190 : std_logic_vector(0 to 0) := (others => '0');
    variable r4189 : std_logic_vector(0 to 0) := (others => '0');
    variable r4188 : std_logic_vector(0 to 0) := (others => '0');
    variable r4187 : std_logic_vector(0 to 0) := (others => '0');
    variable r4186 : std_logic_vector(0 to 0) := (others => '0');
    variable r4185 : std_logic_vector(0 to 0) := (others => '0');
    variable r4184 : std_logic_vector(0 to 0) := (others => '0');
    variable r4183 : std_logic_vector(0 to 0) := (others => '0');
    variable r4182 : std_logic_vector(0 to 0) := (others => '0');
    variable r4181 : std_logic_vector(0 to 0) := (others => '0');
    variable r4180 : std_logic_vector(0 to 0) := (others => '0');
    variable r4179 : std_logic_vector(0 to 0) := (others => '0');
    variable r4178 : std_logic_vector(0 to 0) := (others => '0');
    variable r4177 : std_logic_vector(0 to 0) := (others => '0');
    variable r4176 : std_logic_vector(0 to 0) := (others => '0');
    variable r4175 : std_logic_vector(0 to 0) := (others => '0');
    variable r4174 : std_logic_vector(0 to 0) := (others => '0');
    variable r4173 : std_logic_vector(0 to 0) := (others => '0');
    variable r4172 : std_logic_vector(0 to 0) := (others => '0');
    variable r4171 : std_logic_vector(0 to 0) := (others => '0');
    variable r4170 : std_logic_vector(0 to 0) := (others => '0');
    variable r4169 : std_logic_vector(0 to 0) := (others => '0');
    variable r4168 : std_logic_vector(0 to 0) := (others => '0');
    variable r4167 : std_logic_vector(0 to 0) := (others => '0');
    variable r4166 : std_logic_vector(0 to 0) := (others => '0');
    variable r4165 : std_logic_vector(0 to 0) := (others => '0');
    variable r4164 : std_logic_vector(0 to 0) := (others => '0');
    variable r4163 : std_logic_vector(0 to 0) := (others => '0');
    variable r4162 : std_logic_vector(0 to 0) := (others => '0');
    variable r4161 : std_logic_vector(0 to 0) := (others => '0');
    variable r4160 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r4161 := "0";
    null;
    r4162 := (r4161);
    r4163 := "1";
    null;
    r4164 := (r4163);
    r4165 := "1";
    null;
    r4166 := (r4165);
    r4167 := "0";
    null;
    r4168 := (r4167);
    r4169 := "0";
    null;
    r4170 := (r4169);
    r4171 := "1";
    null;
    r4172 := (r4171);
    r4173 := "0";
    null;
    r4174 := (r4173);
    r4175 := "1";
    null;
    r4176 := (r4175);
    r4177 := "0";
    null;
    r4178 := (r4177);
    r4179 := "0";
    null;
    r4180 := (r4179);
    r4181 := "0";
    null;
    r4182 := (r4181);
    r4183 := "0";
    null;
    r4184 := (r4183);
    r4185 := "1";
    null;
    r4186 := (r4185);
    r4187 := "0";
    null;
    r4188 := (r4187);
    r4189 := "1";
    null;
    r4190 := (r4189);
    r4191 := "0";
    null;
    r4192 := (r4191);
    r4193 := "0";
    null;
    r4194 := (r4193);
    r4195 := "1";
    null;
    r4196 := (r4195);
    r4197 := "1";
    null;
    r4198 := (r4197);
    r4199 := "1";
    null;
    r4200 := (r4199);
    r4201 := "0";
    null;
    r4202 := (r4201);
    r4203 := "0";
    null;
    r4204 := (r4203);
    r4205 := "1";
    null;
    r4206 := (r4205);
    r4207 := "1";
    null;
    r4208 := (r4207);
    r4209 := "0";
    null;
    r4210 := (r4209);
    r4211 := "1";
    null;
    r4212 := (r4211);
    r4213 := "0";
    null;
    r4214 := (r4213);
    r4215 := "1";
    null;
    r4216 := (r4215);
    r4217 := "0";
    null;
    r4218 := (r4217);
    r4219 := "1";
    null;
    r4220 := (r4219);
    r4221 := "0";
    null;
    r4222 := (r4221);
    r4223 := "0";
    null;
    r4224 := (r4223);
    r4160 := (r4162 & r4164 & r4166 & r4168 & r4170 & r4172 & r4174 & r4176 & r4178 & r4180 & r4182 & r4184 & r4186 & r4188 & r4190 & r4192 & r4194 & r4196 & r4198 & r4200 & r4202 & r4204 & r4206 & r4208 & r4210 & r4212 & r4214 & r4216 & r4218 & r4220 & r4222 & r4224);
    return r4160;
  end rewire_MetaprogrammingRW.w650a7354_4159;
  function rewire_MetaprogrammingRW.w53380d13_4090 return std_logic_vector
  is
    variable r4155 : std_logic_vector(0 to 0) := (others => '0');
    variable r4154 : std_logic_vector(0 to 0) := (others => '0');
    variable r4153 : std_logic_vector(0 to 0) := (others => '0');
    variable r4152 : std_logic_vector(0 to 0) := (others => '0');
    variable r4151 : std_logic_vector(0 to 0) := (others => '0');
    variable r4150 : std_logic_vector(0 to 0) := (others => '0');
    variable r4149 : std_logic_vector(0 to 0) := (others => '0');
    variable r4148 : std_logic_vector(0 to 0) := (others => '0');
    variable r4147 : std_logic_vector(0 to 0) := (others => '0');
    variable r4146 : std_logic_vector(0 to 0) := (others => '0');
    variable r4145 : std_logic_vector(0 to 0) := (others => '0');
    variable r4144 : std_logic_vector(0 to 0) := (others => '0');
    variable r4143 : std_logic_vector(0 to 0) := (others => '0');
    variable r4142 : std_logic_vector(0 to 0) := (others => '0');
    variable r4141 : std_logic_vector(0 to 0) := (others => '0');
    variable r4140 : std_logic_vector(0 to 0) := (others => '0');
    variable r4139 : std_logic_vector(0 to 0) := (others => '0');
    variable r4138 : std_logic_vector(0 to 0) := (others => '0');
    variable r4137 : std_logic_vector(0 to 0) := (others => '0');
    variable r4136 : std_logic_vector(0 to 0) := (others => '0');
    variable r4135 : std_logic_vector(0 to 0) := (others => '0');
    variable r4134 : std_logic_vector(0 to 0) := (others => '0');
    variable r4133 : std_logic_vector(0 to 0) := (others => '0');
    variable r4132 : std_logic_vector(0 to 0) := (others => '0');
    variable r4131 : std_logic_vector(0 to 0) := (others => '0');
    variable r4130 : std_logic_vector(0 to 0) := (others => '0');
    variable r4129 : std_logic_vector(0 to 0) := (others => '0');
    variable r4128 : std_logic_vector(0 to 0) := (others => '0');
    variable r4127 : std_logic_vector(0 to 0) := (others => '0');
    variable r4126 : std_logic_vector(0 to 0) := (others => '0');
    variable r4125 : std_logic_vector(0 to 0) := (others => '0');
    variable r4124 : std_logic_vector(0 to 0) := (others => '0');
    variable r4123 : std_logic_vector(0 to 0) := (others => '0');
    variable r4122 : std_logic_vector(0 to 0) := (others => '0');
    variable r4121 : std_logic_vector(0 to 0) := (others => '0');
    variable r4120 : std_logic_vector(0 to 0) := (others => '0');
    variable r4119 : std_logic_vector(0 to 0) := (others => '0');
    variable r4118 : std_logic_vector(0 to 0) := (others => '0');
    variable r4117 : std_logic_vector(0 to 0) := (others => '0');
    variable r4116 : std_logic_vector(0 to 0) := (others => '0');
    variable r4115 : std_logic_vector(0 to 0) := (others => '0');
    variable r4114 : std_logic_vector(0 to 0) := (others => '0');
    variable r4113 : std_logic_vector(0 to 0) := (others => '0');
    variable r4112 : std_logic_vector(0 to 0) := (others => '0');
    variable r4111 : std_logic_vector(0 to 0) := (others => '0');
    variable r4110 : std_logic_vector(0 to 0) := (others => '0');
    variable r4109 : std_logic_vector(0 to 0) := (others => '0');
    variable r4108 : std_logic_vector(0 to 0) := (others => '0');
    variable r4107 : std_logic_vector(0 to 0) := (others => '0');
    variable r4106 : std_logic_vector(0 to 0) := (others => '0');
    variable r4105 : std_logic_vector(0 to 0) := (others => '0');
    variable r4104 : std_logic_vector(0 to 0) := (others => '0');
    variable r4103 : std_logic_vector(0 to 0) := (others => '0');
    variable r4102 : std_logic_vector(0 to 0) := (others => '0');
    variable r4101 : std_logic_vector(0 to 0) := (others => '0');
    variable r4100 : std_logic_vector(0 to 0) := (others => '0');
    variable r4099 : std_logic_vector(0 to 0) := (others => '0');
    variable r4098 : std_logic_vector(0 to 0) := (others => '0');
    variable r4097 : std_logic_vector(0 to 0) := (others => '0');
    variable r4096 : std_logic_vector(0 to 0) := (others => '0');
    variable r4095 : std_logic_vector(0 to 0) := (others => '0');
    variable r4094 : std_logic_vector(0 to 0) := (others => '0');
    variable r4093 : std_logic_vector(0 to 0) := (others => '0');
    variable r4092 : std_logic_vector(0 to 0) := (others => '0');
    variable r4091 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r4092 := "0";
    null;
    r4093 := (r4092);
    r4094 := "1";
    null;
    r4095 := (r4094);
    r4096 := "0";
    null;
    r4097 := (r4096);
    r4098 := "1";
    null;
    r4099 := (r4098);
    r4100 := "0";
    null;
    r4101 := (r4100);
    r4102 := "0";
    null;
    r4103 := (r4102);
    r4104 := "1";
    null;
    r4105 := (r4104);
    r4106 := "1";
    null;
    r4107 := (r4106);
    r4108 := "0";
    null;
    r4109 := (r4108);
    r4110 := "0";
    null;
    r4111 := (r4110);
    r4112 := "1";
    null;
    r4113 := (r4112);
    r4114 := "1";
    null;
    r4115 := (r4114);
    r4116 := "1";
    null;
    r4117 := (r4116);
    r4118 := "0";
    null;
    r4119 := (r4118);
    r4120 := "0";
    null;
    r4121 := (r4120);
    r4122 := "0";
    null;
    r4123 := (r4122);
    r4124 := "0";
    null;
    r4125 := (r4124);
    r4126 := "0";
    null;
    r4127 := (r4126);
    r4128 := "0";
    null;
    r4129 := (r4128);
    r4130 := "0";
    null;
    r4131 := (r4130);
    r4132 := "1";
    null;
    r4133 := (r4132);
    r4134 := "1";
    null;
    r4135 := (r4134);
    r4136 := "0";
    null;
    r4137 := (r4136);
    r4138 := "1";
    null;
    r4139 := (r4138);
    r4140 := "0";
    null;
    r4141 := (r4140);
    r4142 := "0";
    null;
    r4143 := (r4142);
    r4144 := "0";
    null;
    r4145 := (r4144);
    r4146 := "1";
    null;
    r4147 := (r4146);
    r4148 := "0";
    null;
    r4149 := (r4148);
    r4150 := "0";
    null;
    r4151 := (r4150);
    r4152 := "1";
    null;
    r4153 := (r4152);
    r4154 := "1";
    null;
    r4155 := (r4154);
    r4091 := (r4093 & r4095 & r4097 & r4099 & r4101 & r4103 & r4105 & r4107 & r4109 & r4111 & r4113 & r4115 & r4117 & r4119 & r4121 & r4123 & r4125 & r4127 & r4129 & r4131 & r4133 & r4135 & r4137 & r4139 & r4141 & r4143 & r4145 & r4147 & r4149 & r4151 & r4153 & r4155);
    return r4091;
  end rewire_MetaprogrammingRW.w53380d13_4090;
  function rewire_MetaprogrammingRW.w4d2c6dfc_4021 return std_logic_vector
  is
    variable r4086 : std_logic_vector(0 to 0) := (others => '0');
    variable r4085 : std_logic_vector(0 to 0) := (others => '0');
    variable r4084 : std_logic_vector(0 to 0) := (others => '0');
    variable r4083 : std_logic_vector(0 to 0) := (others => '0');
    variable r4082 : std_logic_vector(0 to 0) := (others => '0');
    variable r4081 : std_logic_vector(0 to 0) := (others => '0');
    variable r4080 : std_logic_vector(0 to 0) := (others => '0');
    variable r4079 : std_logic_vector(0 to 0) := (others => '0');
    variable r4078 : std_logic_vector(0 to 0) := (others => '0');
    variable r4077 : std_logic_vector(0 to 0) := (others => '0');
    variable r4076 : std_logic_vector(0 to 0) := (others => '0');
    variable r4075 : std_logic_vector(0 to 0) := (others => '0');
    variable r4074 : std_logic_vector(0 to 0) := (others => '0');
    variable r4073 : std_logic_vector(0 to 0) := (others => '0');
    variable r4072 : std_logic_vector(0 to 0) := (others => '0');
    variable r4071 : std_logic_vector(0 to 0) := (others => '0');
    variable r4070 : std_logic_vector(0 to 0) := (others => '0');
    variable r4069 : std_logic_vector(0 to 0) := (others => '0');
    variable r4068 : std_logic_vector(0 to 0) := (others => '0');
    variable r4067 : std_logic_vector(0 to 0) := (others => '0');
    variable r4066 : std_logic_vector(0 to 0) := (others => '0');
    variable r4065 : std_logic_vector(0 to 0) := (others => '0');
    variable r4064 : std_logic_vector(0 to 0) := (others => '0');
    variable r4063 : std_logic_vector(0 to 0) := (others => '0');
    variable r4062 : std_logic_vector(0 to 0) := (others => '0');
    variable r4061 : std_logic_vector(0 to 0) := (others => '0');
    variable r4060 : std_logic_vector(0 to 0) := (others => '0');
    variable r4059 : std_logic_vector(0 to 0) := (others => '0');
    variable r4058 : std_logic_vector(0 to 0) := (others => '0');
    variable r4057 : std_logic_vector(0 to 0) := (others => '0');
    variable r4056 : std_logic_vector(0 to 0) := (others => '0');
    variable r4055 : std_logic_vector(0 to 0) := (others => '0');
    variable r4054 : std_logic_vector(0 to 0) := (others => '0');
    variable r4053 : std_logic_vector(0 to 0) := (others => '0');
    variable r4052 : std_logic_vector(0 to 0) := (others => '0');
    variable r4051 : std_logic_vector(0 to 0) := (others => '0');
    variable r4050 : std_logic_vector(0 to 0) := (others => '0');
    variable r4049 : std_logic_vector(0 to 0) := (others => '0');
    variable r4048 : std_logic_vector(0 to 0) := (others => '0');
    variable r4047 : std_logic_vector(0 to 0) := (others => '0');
    variable r4046 : std_logic_vector(0 to 0) := (others => '0');
    variable r4045 : std_logic_vector(0 to 0) := (others => '0');
    variable r4044 : std_logic_vector(0 to 0) := (others => '0');
    variable r4043 : std_logic_vector(0 to 0) := (others => '0');
    variable r4042 : std_logic_vector(0 to 0) := (others => '0');
    variable r4041 : std_logic_vector(0 to 0) := (others => '0');
    variable r4040 : std_logic_vector(0 to 0) := (others => '0');
    variable r4039 : std_logic_vector(0 to 0) := (others => '0');
    variable r4038 : std_logic_vector(0 to 0) := (others => '0');
    variable r4037 : std_logic_vector(0 to 0) := (others => '0');
    variable r4036 : std_logic_vector(0 to 0) := (others => '0');
    variable r4035 : std_logic_vector(0 to 0) := (others => '0');
    variable r4034 : std_logic_vector(0 to 0) := (others => '0');
    variable r4033 : std_logic_vector(0 to 0) := (others => '0');
    variable r4032 : std_logic_vector(0 to 0) := (others => '0');
    variable r4031 : std_logic_vector(0 to 0) := (others => '0');
    variable r4030 : std_logic_vector(0 to 0) := (others => '0');
    variable r4029 : std_logic_vector(0 to 0) := (others => '0');
    variable r4028 : std_logic_vector(0 to 0) := (others => '0');
    variable r4027 : std_logic_vector(0 to 0) := (others => '0');
    variable r4026 : std_logic_vector(0 to 0) := (others => '0');
    variable r4025 : std_logic_vector(0 to 0) := (others => '0');
    variable r4024 : std_logic_vector(0 to 0) := (others => '0');
    variable r4023 : std_logic_vector(0 to 0) := (others => '0');
    variable r4022 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r4023 := "0";
    null;
    r4024 := (r4023);
    r4025 := "1";
    null;
    r4026 := (r4025);
    r4027 := "0";
    null;
    r4028 := (r4027);
    r4029 := "0";
    null;
    r4030 := (r4029);
    r4031 := "1";
    null;
    r4032 := (r4031);
    r4033 := "1";
    null;
    r4034 := (r4033);
    r4035 := "0";
    null;
    r4036 := (r4035);
    r4037 := "1";
    null;
    r4038 := (r4037);
    r4039 := "0";
    null;
    r4040 := (r4039);
    r4041 := "0";
    null;
    r4042 := (r4041);
    r4043 := "1";
    null;
    r4044 := (r4043);
    r4045 := "0";
    null;
    r4046 := (r4045);
    r4047 := "1";
    null;
    r4048 := (r4047);
    r4049 := "1";
    null;
    r4050 := (r4049);
    r4051 := "0";
    null;
    r4052 := (r4051);
    r4053 := "0";
    null;
    r4054 := (r4053);
    r4055 := "0";
    null;
    r4056 := (r4055);
    r4057 := "1";
    null;
    r4058 := (r4057);
    r4059 := "1";
    null;
    r4060 := (r4059);
    r4061 := "0";
    null;
    r4062 := (r4061);
    r4063 := "1";
    null;
    r4064 := (r4063);
    r4065 := "1";
    null;
    r4066 := (r4065);
    r4067 := "0";
    null;
    r4068 := (r4067);
    r4069 := "1";
    null;
    r4070 := (r4069);
    r4071 := "1";
    null;
    r4072 := (r4071);
    r4073 := "1";
    null;
    r4074 := (r4073);
    r4075 := "1";
    null;
    r4076 := (r4075);
    r4077 := "1";
    null;
    r4078 := (r4077);
    r4079 := "1";
    null;
    r4080 := (r4079);
    r4081 := "1";
    null;
    r4082 := (r4081);
    r4083 := "0";
    null;
    r4084 := (r4083);
    r4085 := "0";
    null;
    r4086 := (r4085);
    r4022 := (r4024 & r4026 & r4028 & r4030 & r4032 & r4034 & r4036 & r4038 & r4040 & r4042 & r4044 & r4046 & r4048 & r4050 & r4052 & r4054 & r4056 & r4058 & r4060 & r4062 & r4064 & r4066 & r4068 & r4070 & r4072 & r4074 & r4076 & r4078 & r4080 & r4082 & r4084 & r4086);
    return r4022;
  end rewire_MetaprogrammingRW.w4d2c6dfc_4021;
  function rewire_MetaprogrammingRW.w2e1b2138_3952 return std_logic_vector
  is
    variable r4017 : std_logic_vector(0 to 0) := (others => '0');
    variable r4016 : std_logic_vector(0 to 0) := (others => '0');
    variable r4015 : std_logic_vector(0 to 0) := (others => '0');
    variable r4014 : std_logic_vector(0 to 0) := (others => '0');
    variable r4013 : std_logic_vector(0 to 0) := (others => '0');
    variable r4012 : std_logic_vector(0 to 0) := (others => '0');
    variable r4011 : std_logic_vector(0 to 0) := (others => '0');
    variable r4010 : std_logic_vector(0 to 0) := (others => '0');
    variable r4009 : std_logic_vector(0 to 0) := (others => '0');
    variable r4008 : std_logic_vector(0 to 0) := (others => '0');
    variable r4007 : std_logic_vector(0 to 0) := (others => '0');
    variable r4006 : std_logic_vector(0 to 0) := (others => '0');
    variable r4005 : std_logic_vector(0 to 0) := (others => '0');
    variable r4004 : std_logic_vector(0 to 0) := (others => '0');
    variable r4003 : std_logic_vector(0 to 0) := (others => '0');
    variable r4002 : std_logic_vector(0 to 0) := (others => '0');
    variable r4001 : std_logic_vector(0 to 0) := (others => '0');
    variable r4000 : std_logic_vector(0 to 0) := (others => '0');
    variable r3999 : std_logic_vector(0 to 0) := (others => '0');
    variable r3998 : std_logic_vector(0 to 0) := (others => '0');
    variable r3997 : std_logic_vector(0 to 0) := (others => '0');
    variable r3996 : std_logic_vector(0 to 0) := (others => '0');
    variable r3995 : std_logic_vector(0 to 0) := (others => '0');
    variable r3994 : std_logic_vector(0 to 0) := (others => '0');
    variable r3993 : std_logic_vector(0 to 0) := (others => '0');
    variable r3992 : std_logic_vector(0 to 0) := (others => '0');
    variable r3991 : std_logic_vector(0 to 0) := (others => '0');
    variable r3990 : std_logic_vector(0 to 0) := (others => '0');
    variable r3989 : std_logic_vector(0 to 0) := (others => '0');
    variable r3988 : std_logic_vector(0 to 0) := (others => '0');
    variable r3987 : std_logic_vector(0 to 0) := (others => '0');
    variable r3986 : std_logic_vector(0 to 0) := (others => '0');
    variable r3985 : std_logic_vector(0 to 0) := (others => '0');
    variable r3984 : std_logic_vector(0 to 0) := (others => '0');
    variable r3983 : std_logic_vector(0 to 0) := (others => '0');
    variable r3982 : std_logic_vector(0 to 0) := (others => '0');
    variable r3981 : std_logic_vector(0 to 0) := (others => '0');
    variable r3980 : std_logic_vector(0 to 0) := (others => '0');
    variable r3979 : std_logic_vector(0 to 0) := (others => '0');
    variable r3978 : std_logic_vector(0 to 0) := (others => '0');
    variable r3977 : std_logic_vector(0 to 0) := (others => '0');
    variable r3976 : std_logic_vector(0 to 0) := (others => '0');
    variable r3975 : std_logic_vector(0 to 0) := (others => '0');
    variable r3974 : std_logic_vector(0 to 0) := (others => '0');
    variable r3973 : std_logic_vector(0 to 0) := (others => '0');
    variable r3972 : std_logic_vector(0 to 0) := (others => '0');
    variable r3971 : std_logic_vector(0 to 0) := (others => '0');
    variable r3970 : std_logic_vector(0 to 0) := (others => '0');
    variable r3969 : std_logic_vector(0 to 0) := (others => '0');
    variable r3968 : std_logic_vector(0 to 0) := (others => '0');
    variable r3967 : std_logic_vector(0 to 0) := (others => '0');
    variable r3966 : std_logic_vector(0 to 0) := (others => '0');
    variable r3965 : std_logic_vector(0 to 0) := (others => '0');
    variable r3964 : std_logic_vector(0 to 0) := (others => '0');
    variable r3963 : std_logic_vector(0 to 0) := (others => '0');
    variable r3962 : std_logic_vector(0 to 0) := (others => '0');
    variable r3961 : std_logic_vector(0 to 0) := (others => '0');
    variable r3960 : std_logic_vector(0 to 0) := (others => '0');
    variable r3959 : std_logic_vector(0 to 0) := (others => '0');
    variable r3958 : std_logic_vector(0 to 0) := (others => '0');
    variable r3957 : std_logic_vector(0 to 0) := (others => '0');
    variable r3956 : std_logic_vector(0 to 0) := (others => '0');
    variable r3955 : std_logic_vector(0 to 0) := (others => '0');
    variable r3954 : std_logic_vector(0 to 0) := (others => '0');
    variable r3953 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r3954 := "0";
    null;
    r3955 := (r3954);
    r3956 := "0";
    null;
    r3957 := (r3956);
    r3958 := "1";
    null;
    r3959 := (r3958);
    r3960 := "0";
    null;
    r3961 := (r3960);
    r3962 := "1";
    null;
    r3963 := (r3962);
    r3964 := "1";
    null;
    r3965 := (r3964);
    r3966 := "1";
    null;
    r3967 := (r3966);
    r3968 := "0";
    null;
    r3969 := (r3968);
    r3970 := "0";
    null;
    r3971 := (r3970);
    r3972 := "0";
    null;
    r3973 := (r3972);
    r3974 := "0";
    null;
    r3975 := (r3974);
    r3976 := "1";
    null;
    r3977 := (r3976);
    r3978 := "1";
    null;
    r3979 := (r3978);
    r3980 := "0";
    null;
    r3981 := (r3980);
    r3982 := "1";
    null;
    r3983 := (r3982);
    r3984 := "1";
    null;
    r3985 := (r3984);
    r3986 := "0";
    null;
    r3987 := (r3986);
    r3988 := "0";
    null;
    r3989 := (r3988);
    r3990 := "1";
    null;
    r3991 := (r3990);
    r3992 := "0";
    null;
    r3993 := (r3992);
    r3994 := "0";
    null;
    r3995 := (r3994);
    r3996 := "0";
    null;
    r3997 := (r3996);
    r3998 := "0";
    null;
    r3999 := (r3998);
    r4000 := "1";
    null;
    r4001 := (r4000);
    r4002 := "0";
    null;
    r4003 := (r4002);
    r4004 := "0";
    null;
    r4005 := (r4004);
    r4006 := "1";
    null;
    r4007 := (r4006);
    r4008 := "1";
    null;
    r4009 := (r4008);
    r4010 := "1";
    null;
    r4011 := (r4010);
    r4012 := "0";
    null;
    r4013 := (r4012);
    r4014 := "0";
    null;
    r4015 := (r4014);
    r4016 := "0";
    null;
    r4017 := (r4016);
    r3953 := (r3955 & r3957 & r3959 & r3961 & r3963 & r3965 & r3967 & r3969 & r3971 & r3973 & r3975 & r3977 & r3979 & r3981 & r3983 & r3985 & r3987 & r3989 & r3991 & r3993 & r3995 & r3997 & r3999 & r4001 & r4003 & r4005 & r4007 & r4009 & r4011 & r4013 & r4015 & r4017);
    return r3953;
  end rewire_MetaprogrammingRW.w2e1b2138_3952;
  function rewire_MetaprogrammingRW.w27b70a85_3883 return std_logic_vector
  is
    variable r3948 : std_logic_vector(0 to 0) := (others => '0');
    variable r3947 : std_logic_vector(0 to 0) := (others => '0');
    variable r3946 : std_logic_vector(0 to 0) := (others => '0');
    variable r3945 : std_logic_vector(0 to 0) := (others => '0');
    variable r3944 : std_logic_vector(0 to 0) := (others => '0');
    variable r3943 : std_logic_vector(0 to 0) := (others => '0');
    variable r3942 : std_logic_vector(0 to 0) := (others => '0');
    variable r3941 : std_logic_vector(0 to 0) := (others => '0');
    variable r3940 : std_logic_vector(0 to 0) := (others => '0');
    variable r3939 : std_logic_vector(0 to 0) := (others => '0');
    variable r3938 : std_logic_vector(0 to 0) := (others => '0');
    variable r3937 : std_logic_vector(0 to 0) := (others => '0');
    variable r3936 : std_logic_vector(0 to 0) := (others => '0');
    variable r3935 : std_logic_vector(0 to 0) := (others => '0');
    variable r3934 : std_logic_vector(0 to 0) := (others => '0');
    variable r3933 : std_logic_vector(0 to 0) := (others => '0');
    variable r3932 : std_logic_vector(0 to 0) := (others => '0');
    variable r3931 : std_logic_vector(0 to 0) := (others => '0');
    variable r3930 : std_logic_vector(0 to 0) := (others => '0');
    variable r3929 : std_logic_vector(0 to 0) := (others => '0');
    variable r3928 : std_logic_vector(0 to 0) := (others => '0');
    variable r3927 : std_logic_vector(0 to 0) := (others => '0');
    variable r3926 : std_logic_vector(0 to 0) := (others => '0');
    variable r3925 : std_logic_vector(0 to 0) := (others => '0');
    variable r3924 : std_logic_vector(0 to 0) := (others => '0');
    variable r3923 : std_logic_vector(0 to 0) := (others => '0');
    variable r3922 : std_logic_vector(0 to 0) := (others => '0');
    variable r3921 : std_logic_vector(0 to 0) := (others => '0');
    variable r3920 : std_logic_vector(0 to 0) := (others => '0');
    variable r3919 : std_logic_vector(0 to 0) := (others => '0');
    variable r3918 : std_logic_vector(0 to 0) := (others => '0');
    variable r3917 : std_logic_vector(0 to 0) := (others => '0');
    variable r3916 : std_logic_vector(0 to 0) := (others => '0');
    variable r3915 : std_logic_vector(0 to 0) := (others => '0');
    variable r3914 : std_logic_vector(0 to 0) := (others => '0');
    variable r3913 : std_logic_vector(0 to 0) := (others => '0');
    variable r3912 : std_logic_vector(0 to 0) := (others => '0');
    variable r3911 : std_logic_vector(0 to 0) := (others => '0');
    variable r3910 : std_logic_vector(0 to 0) := (others => '0');
    variable r3909 : std_logic_vector(0 to 0) := (others => '0');
    variable r3908 : std_logic_vector(0 to 0) := (others => '0');
    variable r3907 : std_logic_vector(0 to 0) := (others => '0');
    variable r3906 : std_logic_vector(0 to 0) := (others => '0');
    variable r3905 : std_logic_vector(0 to 0) := (others => '0');
    variable r3904 : std_logic_vector(0 to 0) := (others => '0');
    variable r3903 : std_logic_vector(0 to 0) := (others => '0');
    variable r3902 : std_logic_vector(0 to 0) := (others => '0');
    variable r3901 : std_logic_vector(0 to 0) := (others => '0');
    variable r3900 : std_logic_vector(0 to 0) := (others => '0');
    variable r3899 : std_logic_vector(0 to 0) := (others => '0');
    variable r3898 : std_logic_vector(0 to 0) := (others => '0');
    variable r3897 : std_logic_vector(0 to 0) := (others => '0');
    variable r3896 : std_logic_vector(0 to 0) := (others => '0');
    variable r3895 : std_logic_vector(0 to 0) := (others => '0');
    variable r3894 : std_logic_vector(0 to 0) := (others => '0');
    variable r3893 : std_logic_vector(0 to 0) := (others => '0');
    variable r3892 : std_logic_vector(0 to 0) := (others => '0');
    variable r3891 : std_logic_vector(0 to 0) := (others => '0');
    variable r3890 : std_logic_vector(0 to 0) := (others => '0');
    variable r3889 : std_logic_vector(0 to 0) := (others => '0');
    variable r3888 : std_logic_vector(0 to 0) := (others => '0');
    variable r3887 : std_logic_vector(0 to 0) := (others => '0');
    variable r3886 : std_logic_vector(0 to 0) := (others => '0');
    variable r3885 : std_logic_vector(0 to 0) := (others => '0');
    variable r3884 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r3885 := "0";
    null;
    r3886 := (r3885);
    r3887 := "0";
    null;
    r3888 := (r3887);
    r3889 := "1";
    null;
    r3890 := (r3889);
    r3891 := "0";
    null;
    r3892 := (r3891);
    r3893 := "0";
    null;
    r3894 := (r3893);
    r3895 := "1";
    null;
    r3896 := (r3895);
    r3897 := "1";
    null;
    r3898 := (r3897);
    r3899 := "1";
    null;
    r3900 := (r3899);
    r3901 := "1";
    null;
    r3902 := (r3901);
    r3903 := "0";
    null;
    r3904 := (r3903);
    r3905 := "1";
    null;
    r3906 := (r3905);
    r3907 := "1";
    null;
    r3908 := (r3907);
    r3909 := "0";
    null;
    r3910 := (r3909);
    r3911 := "1";
    null;
    r3912 := (r3911);
    r3913 := "1";
    null;
    r3914 := (r3913);
    r3915 := "1";
    null;
    r3916 := (r3915);
    r3917 := "0";
    null;
    r3918 := (r3917);
    r3919 := "0";
    null;
    r3920 := (r3919);
    r3921 := "0";
    null;
    r3922 := (r3921);
    r3923 := "0";
    null;
    r3924 := (r3923);
    r3925 := "1";
    null;
    r3926 := (r3925);
    r3927 := "0";
    null;
    r3928 := (r3927);
    r3929 := "1";
    null;
    r3930 := (r3929);
    r3931 := "0";
    null;
    r3932 := (r3931);
    r3933 := "1";
    null;
    r3934 := (r3933);
    r3935 := "0";
    null;
    r3936 := (r3935);
    r3937 := "0";
    null;
    r3938 := (r3937);
    r3939 := "0";
    null;
    r3940 := (r3939);
    r3941 := "0";
    null;
    r3942 := (r3941);
    r3943 := "1";
    null;
    r3944 := (r3943);
    r3945 := "0";
    null;
    r3946 := (r3945);
    r3947 := "1";
    null;
    r3948 := (r3947);
    r3884 := (r3886 & r3888 & r3890 & r3892 & r3894 & r3896 & r3898 & r3900 & r3902 & r3904 & r3906 & r3908 & r3910 & r3912 & r3914 & r3916 & r3918 & r3920 & r3922 & r3924 & r3926 & r3928 & r3930 & r3932 & r3934 & r3936 & r3938 & r3940 & r3942 & r3944 & r3946 & r3948);
    return r3884;
  end rewire_MetaprogrammingRW.w27b70a85_3883;
  function rewire_MetaprogrammingRW.w14292967_3814 return std_logic_vector
  is
    variable r3879 : std_logic_vector(0 to 0) := (others => '0');
    variable r3878 : std_logic_vector(0 to 0) := (others => '0');
    variable r3877 : std_logic_vector(0 to 0) := (others => '0');
    variable r3876 : std_logic_vector(0 to 0) := (others => '0');
    variable r3875 : std_logic_vector(0 to 0) := (others => '0');
    variable r3874 : std_logic_vector(0 to 0) := (others => '0');
    variable r3873 : std_logic_vector(0 to 0) := (others => '0');
    variable r3872 : std_logic_vector(0 to 0) := (others => '0');
    variable r3871 : std_logic_vector(0 to 0) := (others => '0');
    variable r3870 : std_logic_vector(0 to 0) := (others => '0');
    variable r3869 : std_logic_vector(0 to 0) := (others => '0');
    variable r3868 : std_logic_vector(0 to 0) := (others => '0');
    variable r3867 : std_logic_vector(0 to 0) := (others => '0');
    variable r3866 : std_logic_vector(0 to 0) := (others => '0');
    variable r3865 : std_logic_vector(0 to 0) := (others => '0');
    variable r3864 : std_logic_vector(0 to 0) := (others => '0');
    variable r3863 : std_logic_vector(0 to 0) := (others => '0');
    variable r3862 : std_logic_vector(0 to 0) := (others => '0');
    variable r3861 : std_logic_vector(0 to 0) := (others => '0');
    variable r3860 : std_logic_vector(0 to 0) := (others => '0');
    variable r3859 : std_logic_vector(0 to 0) := (others => '0');
    variable r3858 : std_logic_vector(0 to 0) := (others => '0');
    variable r3857 : std_logic_vector(0 to 0) := (others => '0');
    variable r3856 : std_logic_vector(0 to 0) := (others => '0');
    variable r3855 : std_logic_vector(0 to 0) := (others => '0');
    variable r3854 : std_logic_vector(0 to 0) := (others => '0');
    variable r3853 : std_logic_vector(0 to 0) := (others => '0');
    variable r3852 : std_logic_vector(0 to 0) := (others => '0');
    variable r3851 : std_logic_vector(0 to 0) := (others => '0');
    variable r3850 : std_logic_vector(0 to 0) := (others => '0');
    variable r3849 : std_logic_vector(0 to 0) := (others => '0');
    variable r3848 : std_logic_vector(0 to 0) := (others => '0');
    variable r3847 : std_logic_vector(0 to 0) := (others => '0');
    variable r3846 : std_logic_vector(0 to 0) := (others => '0');
    variable r3845 : std_logic_vector(0 to 0) := (others => '0');
    variable r3844 : std_logic_vector(0 to 0) := (others => '0');
    variable r3843 : std_logic_vector(0 to 0) := (others => '0');
    variable r3842 : std_logic_vector(0 to 0) := (others => '0');
    variable r3841 : std_logic_vector(0 to 0) := (others => '0');
    variable r3840 : std_logic_vector(0 to 0) := (others => '0');
    variable r3839 : std_logic_vector(0 to 0) := (others => '0');
    variable r3838 : std_logic_vector(0 to 0) := (others => '0');
    variable r3837 : std_logic_vector(0 to 0) := (others => '0');
    variable r3836 : std_logic_vector(0 to 0) := (others => '0');
    variable r3835 : std_logic_vector(0 to 0) := (others => '0');
    variable r3834 : std_logic_vector(0 to 0) := (others => '0');
    variable r3833 : std_logic_vector(0 to 0) := (others => '0');
    variable r3832 : std_logic_vector(0 to 0) := (others => '0');
    variable r3831 : std_logic_vector(0 to 0) := (others => '0');
    variable r3830 : std_logic_vector(0 to 0) := (others => '0');
    variable r3829 : std_logic_vector(0 to 0) := (others => '0');
    variable r3828 : std_logic_vector(0 to 0) := (others => '0');
    variable r3827 : std_logic_vector(0 to 0) := (others => '0');
    variable r3826 : std_logic_vector(0 to 0) := (others => '0');
    variable r3825 : std_logic_vector(0 to 0) := (others => '0');
    variable r3824 : std_logic_vector(0 to 0) := (others => '0');
    variable r3823 : std_logic_vector(0 to 0) := (others => '0');
    variable r3822 : std_logic_vector(0 to 0) := (others => '0');
    variable r3821 : std_logic_vector(0 to 0) := (others => '0');
    variable r3820 : std_logic_vector(0 to 0) := (others => '0');
    variable r3819 : std_logic_vector(0 to 0) := (others => '0');
    variable r3818 : std_logic_vector(0 to 0) := (others => '0');
    variable r3817 : std_logic_vector(0 to 0) := (others => '0');
    variable r3816 : std_logic_vector(0 to 0) := (others => '0');
    variable r3815 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r3816 := "0";
    null;
    r3817 := (r3816);
    r3818 := "0";
    null;
    r3819 := (r3818);
    r3820 := "0";
    null;
    r3821 := (r3820);
    r3822 := "1";
    null;
    r3823 := (r3822);
    r3824 := "0";
    null;
    r3825 := (r3824);
    r3826 := "1";
    null;
    r3827 := (r3826);
    r3828 := "0";
    null;
    r3829 := (r3828);
    r3830 := "0";
    null;
    r3831 := (r3830);
    r3832 := "0";
    null;
    r3833 := (r3832);
    r3834 := "0";
    null;
    r3835 := (r3834);
    r3836 := "1";
    null;
    r3837 := (r3836);
    r3838 := "0";
    null;
    r3839 := (r3838);
    r3840 := "1";
    null;
    r3841 := (r3840);
    r3842 := "0";
    null;
    r3843 := (r3842);
    r3844 := "0";
    null;
    r3845 := (r3844);
    r3846 := "1";
    null;
    r3847 := (r3846);
    r3848 := "0";
    null;
    r3849 := (r3848);
    r3850 := "0";
    null;
    r3851 := (r3850);
    r3852 := "1";
    null;
    r3853 := (r3852);
    r3854 := "0";
    null;
    r3855 := (r3854);
    r3856 := "1";
    null;
    r3857 := (r3856);
    r3858 := "0";
    null;
    r3859 := (r3858);
    r3860 := "0";
    null;
    r3861 := (r3860);
    r3862 := "1";
    null;
    r3863 := (r3862);
    r3864 := "0";
    null;
    r3865 := (r3864);
    r3866 := "1";
    null;
    r3867 := (r3866);
    r3868 := "1";
    null;
    r3869 := (r3868);
    r3870 := "0";
    null;
    r3871 := (r3870);
    r3872 := "0";
    null;
    r3873 := (r3872);
    r3874 := "1";
    null;
    r3875 := (r3874);
    r3876 := "1";
    null;
    r3877 := (r3876);
    r3878 := "1";
    null;
    r3879 := (r3878);
    r3815 := (r3817 & r3819 & r3821 & r3823 & r3825 & r3827 & r3829 & r3831 & r3833 & r3835 & r3837 & r3839 & r3841 & r3843 & r3845 & r3847 & r3849 & r3851 & r3853 & r3855 & r3857 & r3859 & r3861 & r3863 & r3865 & r3867 & r3869 & r3871 & r3873 & r3875 & r3877 & r3879);
    return r3815;
  end rewire_MetaprogrammingRW.w14292967_3814;
  function rewire_MetaprogrammingRW.w06ca6351_3745 return std_logic_vector
  is
    variable r3810 : std_logic_vector(0 to 0) := (others => '0');
    variable r3809 : std_logic_vector(0 to 0) := (others => '0');
    variable r3808 : std_logic_vector(0 to 0) := (others => '0');
    variable r3807 : std_logic_vector(0 to 0) := (others => '0');
    variable r3806 : std_logic_vector(0 to 0) := (others => '0');
    variable r3805 : std_logic_vector(0 to 0) := (others => '0');
    variable r3804 : std_logic_vector(0 to 0) := (others => '0');
    variable r3803 : std_logic_vector(0 to 0) := (others => '0');
    variable r3802 : std_logic_vector(0 to 0) := (others => '0');
    variable r3801 : std_logic_vector(0 to 0) := (others => '0');
    variable r3800 : std_logic_vector(0 to 0) := (others => '0');
    variable r3799 : std_logic_vector(0 to 0) := (others => '0');
    variable r3798 : std_logic_vector(0 to 0) := (others => '0');
    variable r3797 : std_logic_vector(0 to 0) := (others => '0');
    variable r3796 : std_logic_vector(0 to 0) := (others => '0');
    variable r3795 : std_logic_vector(0 to 0) := (others => '0');
    variable r3794 : std_logic_vector(0 to 0) := (others => '0');
    variable r3793 : std_logic_vector(0 to 0) := (others => '0');
    variable r3792 : std_logic_vector(0 to 0) := (others => '0');
    variable r3791 : std_logic_vector(0 to 0) := (others => '0');
    variable r3790 : std_logic_vector(0 to 0) := (others => '0');
    variable r3789 : std_logic_vector(0 to 0) := (others => '0');
    variable r3788 : std_logic_vector(0 to 0) := (others => '0');
    variable r3787 : std_logic_vector(0 to 0) := (others => '0');
    variable r3786 : std_logic_vector(0 to 0) := (others => '0');
    variable r3785 : std_logic_vector(0 to 0) := (others => '0');
    variable r3784 : std_logic_vector(0 to 0) := (others => '0');
    variable r3783 : std_logic_vector(0 to 0) := (others => '0');
    variable r3782 : std_logic_vector(0 to 0) := (others => '0');
    variable r3781 : std_logic_vector(0 to 0) := (others => '0');
    variable r3780 : std_logic_vector(0 to 0) := (others => '0');
    variable r3779 : std_logic_vector(0 to 0) := (others => '0');
    variable r3778 : std_logic_vector(0 to 0) := (others => '0');
    variable r3777 : std_logic_vector(0 to 0) := (others => '0');
    variable r3776 : std_logic_vector(0 to 0) := (others => '0');
    variable r3775 : std_logic_vector(0 to 0) := (others => '0');
    variable r3774 : std_logic_vector(0 to 0) := (others => '0');
    variable r3773 : std_logic_vector(0 to 0) := (others => '0');
    variable r3772 : std_logic_vector(0 to 0) := (others => '0');
    variable r3771 : std_logic_vector(0 to 0) := (others => '0');
    variable r3770 : std_logic_vector(0 to 0) := (others => '0');
    variable r3769 : std_logic_vector(0 to 0) := (others => '0');
    variable r3768 : std_logic_vector(0 to 0) := (others => '0');
    variable r3767 : std_logic_vector(0 to 0) := (others => '0');
    variable r3766 : std_logic_vector(0 to 0) := (others => '0');
    variable r3765 : std_logic_vector(0 to 0) := (others => '0');
    variable r3764 : std_logic_vector(0 to 0) := (others => '0');
    variable r3763 : std_logic_vector(0 to 0) := (others => '0');
    variable r3762 : std_logic_vector(0 to 0) := (others => '0');
    variable r3761 : std_logic_vector(0 to 0) := (others => '0');
    variable r3760 : std_logic_vector(0 to 0) := (others => '0');
    variable r3759 : std_logic_vector(0 to 0) := (others => '0');
    variable r3758 : std_logic_vector(0 to 0) := (others => '0');
    variable r3757 : std_logic_vector(0 to 0) := (others => '0');
    variable r3756 : std_logic_vector(0 to 0) := (others => '0');
    variable r3755 : std_logic_vector(0 to 0) := (others => '0');
    variable r3754 : std_logic_vector(0 to 0) := (others => '0');
    variable r3753 : std_logic_vector(0 to 0) := (others => '0');
    variable r3752 : std_logic_vector(0 to 0) := (others => '0');
    variable r3751 : std_logic_vector(0 to 0) := (others => '0');
    variable r3750 : std_logic_vector(0 to 0) := (others => '0');
    variable r3749 : std_logic_vector(0 to 0) := (others => '0');
    variable r3748 : std_logic_vector(0 to 0) := (others => '0');
    variable r3747 : std_logic_vector(0 to 0) := (others => '0');
    variable r3746 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r3747 := "0";
    null;
    r3748 := (r3747);
    r3749 := "0";
    null;
    r3750 := (r3749);
    r3751 := "0";
    null;
    r3752 := (r3751);
    r3753 := "0";
    null;
    r3754 := (r3753);
    r3755 := "0";
    null;
    r3756 := (r3755);
    r3757 := "1";
    null;
    r3758 := (r3757);
    r3759 := "1";
    null;
    r3760 := (r3759);
    r3761 := "0";
    null;
    r3762 := (r3761);
    r3763 := "1";
    null;
    r3764 := (r3763);
    r3765 := "1";
    null;
    r3766 := (r3765);
    r3767 := "0";
    null;
    r3768 := (r3767);
    r3769 := "0";
    null;
    r3770 := (r3769);
    r3771 := "1";
    null;
    r3772 := (r3771);
    r3773 := "0";
    null;
    r3774 := (r3773);
    r3775 := "1";
    null;
    r3776 := (r3775);
    r3777 := "0";
    null;
    r3778 := (r3777);
    r3779 := "0";
    null;
    r3780 := (r3779);
    r3781 := "1";
    null;
    r3782 := (r3781);
    r3783 := "1";
    null;
    r3784 := (r3783);
    r3785 := "0";
    null;
    r3786 := (r3785);
    r3787 := "0";
    null;
    r3788 := (r3787);
    r3789 := "0";
    null;
    r3790 := (r3789);
    r3791 := "1";
    null;
    r3792 := (r3791);
    r3793 := "1";
    null;
    r3794 := (r3793);
    r3795 := "0";
    null;
    r3796 := (r3795);
    r3797 := "1";
    null;
    r3798 := (r3797);
    r3799 := "0";
    null;
    r3800 := (r3799);
    r3801 := "1";
    null;
    r3802 := (r3801);
    r3803 := "0";
    null;
    r3804 := (r3803);
    r3805 := "0";
    null;
    r3806 := (r3805);
    r3807 := "0";
    null;
    r3808 := (r3807);
    r3809 := "1";
    null;
    r3810 := (r3809);
    r3746 := (r3748 & r3750 & r3752 & r3754 & r3756 & r3758 & r3760 & r3762 & r3764 & r3766 & r3768 & r3770 & r3772 & r3774 & r3776 & r3778 & r3780 & r3782 & r3784 & r3786 & r3788 & r3790 & r3792 & r3794 & r3796 & r3798 & r3800 & r3802 & r3804 & r3806 & r3808 & r3810);
    return r3746;
  end rewire_MetaprogrammingRW.w06ca6351_3745;
  function rewire_MetaprogrammingRW.wd5a79147_3676 return std_logic_vector
  is
    variable r3741 : std_logic_vector(0 to 0) := (others => '0');
    variable r3740 : std_logic_vector(0 to 0) := (others => '0');
    variable r3739 : std_logic_vector(0 to 0) := (others => '0');
    variable r3738 : std_logic_vector(0 to 0) := (others => '0');
    variable r3737 : std_logic_vector(0 to 0) := (others => '0');
    variable r3736 : std_logic_vector(0 to 0) := (others => '0');
    variable r3735 : std_logic_vector(0 to 0) := (others => '0');
    variable r3734 : std_logic_vector(0 to 0) := (others => '0');
    variable r3733 : std_logic_vector(0 to 0) := (others => '0');
    variable r3732 : std_logic_vector(0 to 0) := (others => '0');
    variable r3731 : std_logic_vector(0 to 0) := (others => '0');
    variable r3730 : std_logic_vector(0 to 0) := (others => '0');
    variable r3729 : std_logic_vector(0 to 0) := (others => '0');
    variable r3728 : std_logic_vector(0 to 0) := (others => '0');
    variable r3727 : std_logic_vector(0 to 0) := (others => '0');
    variable r3726 : std_logic_vector(0 to 0) := (others => '0');
    variable r3725 : std_logic_vector(0 to 0) := (others => '0');
    variable r3724 : std_logic_vector(0 to 0) := (others => '0');
    variable r3723 : std_logic_vector(0 to 0) := (others => '0');
    variable r3722 : std_logic_vector(0 to 0) := (others => '0');
    variable r3721 : std_logic_vector(0 to 0) := (others => '0');
    variable r3720 : std_logic_vector(0 to 0) := (others => '0');
    variable r3719 : std_logic_vector(0 to 0) := (others => '0');
    variable r3718 : std_logic_vector(0 to 0) := (others => '0');
    variable r3717 : std_logic_vector(0 to 0) := (others => '0');
    variable r3716 : std_logic_vector(0 to 0) := (others => '0');
    variable r3715 : std_logic_vector(0 to 0) := (others => '0');
    variable r3714 : std_logic_vector(0 to 0) := (others => '0');
    variable r3713 : std_logic_vector(0 to 0) := (others => '0');
    variable r3712 : std_logic_vector(0 to 0) := (others => '0');
    variable r3711 : std_logic_vector(0 to 0) := (others => '0');
    variable r3710 : std_logic_vector(0 to 0) := (others => '0');
    variable r3709 : std_logic_vector(0 to 0) := (others => '0');
    variable r3708 : std_logic_vector(0 to 0) := (others => '0');
    variable r3707 : std_logic_vector(0 to 0) := (others => '0');
    variable r3706 : std_logic_vector(0 to 0) := (others => '0');
    variable r3705 : std_logic_vector(0 to 0) := (others => '0');
    variable r3704 : std_logic_vector(0 to 0) := (others => '0');
    variable r3703 : std_logic_vector(0 to 0) := (others => '0');
    variable r3702 : std_logic_vector(0 to 0) := (others => '0');
    variable r3701 : std_logic_vector(0 to 0) := (others => '0');
    variable r3700 : std_logic_vector(0 to 0) := (others => '0');
    variable r3699 : std_logic_vector(0 to 0) := (others => '0');
    variable r3698 : std_logic_vector(0 to 0) := (others => '0');
    variable r3697 : std_logic_vector(0 to 0) := (others => '0');
    variable r3696 : std_logic_vector(0 to 0) := (others => '0');
    variable r3695 : std_logic_vector(0 to 0) := (others => '0');
    variable r3694 : std_logic_vector(0 to 0) := (others => '0');
    variable r3693 : std_logic_vector(0 to 0) := (others => '0');
    variable r3692 : std_logic_vector(0 to 0) := (others => '0');
    variable r3691 : std_logic_vector(0 to 0) := (others => '0');
    variable r3690 : std_logic_vector(0 to 0) := (others => '0');
    variable r3689 : std_logic_vector(0 to 0) := (others => '0');
    variable r3688 : std_logic_vector(0 to 0) := (others => '0');
    variable r3687 : std_logic_vector(0 to 0) := (others => '0');
    variable r3686 : std_logic_vector(0 to 0) := (others => '0');
    variable r3685 : std_logic_vector(0 to 0) := (others => '0');
    variable r3684 : std_logic_vector(0 to 0) := (others => '0');
    variable r3683 : std_logic_vector(0 to 0) := (others => '0');
    variable r3682 : std_logic_vector(0 to 0) := (others => '0');
    variable r3681 : std_logic_vector(0 to 0) := (others => '0');
    variable r3680 : std_logic_vector(0 to 0) := (others => '0');
    variable r3679 : std_logic_vector(0 to 0) := (others => '0');
    variable r3678 : std_logic_vector(0 to 0) := (others => '0');
    variable r3677 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r3678 := "1";
    null;
    r3679 := (r3678);
    r3680 := "1";
    null;
    r3681 := (r3680);
    r3682 := "0";
    null;
    r3683 := (r3682);
    r3684 := "1";
    null;
    r3685 := (r3684);
    r3686 := "0";
    null;
    r3687 := (r3686);
    r3688 := "1";
    null;
    r3689 := (r3688);
    r3690 := "0";
    null;
    r3691 := (r3690);
    r3692 := "1";
    null;
    r3693 := (r3692);
    r3694 := "1";
    null;
    r3695 := (r3694);
    r3696 := "0";
    null;
    r3697 := (r3696);
    r3698 := "1";
    null;
    r3699 := (r3698);
    r3700 := "0";
    null;
    r3701 := (r3700);
    r3702 := "0";
    null;
    r3703 := (r3702);
    r3704 := "1";
    null;
    r3705 := (r3704);
    r3706 := "1";
    null;
    r3707 := (r3706);
    r3708 := "1";
    null;
    r3709 := (r3708);
    r3710 := "1";
    null;
    r3711 := (r3710);
    r3712 := "0";
    null;
    r3713 := (r3712);
    r3714 := "0";
    null;
    r3715 := (r3714);
    r3716 := "1";
    null;
    r3717 := (r3716);
    r3718 := "0";
    null;
    r3719 := (r3718);
    r3720 := "0";
    null;
    r3721 := (r3720);
    r3722 := "0";
    null;
    r3723 := (r3722);
    r3724 := "1";
    null;
    r3725 := (r3724);
    r3726 := "0";
    null;
    r3727 := (r3726);
    r3728 := "1";
    null;
    r3729 := (r3728);
    r3730 := "0";
    null;
    r3731 := (r3730);
    r3732 := "0";
    null;
    r3733 := (r3732);
    r3734 := "0";
    null;
    r3735 := (r3734);
    r3736 := "1";
    null;
    r3737 := (r3736);
    r3738 := "1";
    null;
    r3739 := (r3738);
    r3740 := "1";
    null;
    r3741 := (r3740);
    r3677 := (r3679 & r3681 & r3683 & r3685 & r3687 & r3689 & r3691 & r3693 & r3695 & r3697 & r3699 & r3701 & r3703 & r3705 & r3707 & r3709 & r3711 & r3713 & r3715 & r3717 & r3719 & r3721 & r3723 & r3725 & r3727 & r3729 & r3731 & r3733 & r3735 & r3737 & r3739 & r3741);
    return r3677;
  end rewire_MetaprogrammingRW.wd5a79147_3676;
  function rewire_MetaprogrammingRW.wc6e00bf3_3607 return std_logic_vector
  is
    variable r3672 : std_logic_vector(0 to 0) := (others => '0');
    variable r3671 : std_logic_vector(0 to 0) := (others => '0');
    variable r3670 : std_logic_vector(0 to 0) := (others => '0');
    variable r3669 : std_logic_vector(0 to 0) := (others => '0');
    variable r3668 : std_logic_vector(0 to 0) := (others => '0');
    variable r3667 : std_logic_vector(0 to 0) := (others => '0');
    variable r3666 : std_logic_vector(0 to 0) := (others => '0');
    variable r3665 : std_logic_vector(0 to 0) := (others => '0');
    variable r3664 : std_logic_vector(0 to 0) := (others => '0');
    variable r3663 : std_logic_vector(0 to 0) := (others => '0');
    variable r3662 : std_logic_vector(0 to 0) := (others => '0');
    variable r3661 : std_logic_vector(0 to 0) := (others => '0');
    variable r3660 : std_logic_vector(0 to 0) := (others => '0');
    variable r3659 : std_logic_vector(0 to 0) := (others => '0');
    variable r3658 : std_logic_vector(0 to 0) := (others => '0');
    variable r3657 : std_logic_vector(0 to 0) := (others => '0');
    variable r3656 : std_logic_vector(0 to 0) := (others => '0');
    variable r3655 : std_logic_vector(0 to 0) := (others => '0');
    variable r3654 : std_logic_vector(0 to 0) := (others => '0');
    variable r3653 : std_logic_vector(0 to 0) := (others => '0');
    variable r3652 : std_logic_vector(0 to 0) := (others => '0');
    variable r3651 : std_logic_vector(0 to 0) := (others => '0');
    variable r3650 : std_logic_vector(0 to 0) := (others => '0');
    variable r3649 : std_logic_vector(0 to 0) := (others => '0');
    variable r3648 : std_logic_vector(0 to 0) := (others => '0');
    variable r3647 : std_logic_vector(0 to 0) := (others => '0');
    variable r3646 : std_logic_vector(0 to 0) := (others => '0');
    variable r3645 : std_logic_vector(0 to 0) := (others => '0');
    variable r3644 : std_logic_vector(0 to 0) := (others => '0');
    variable r3643 : std_logic_vector(0 to 0) := (others => '0');
    variable r3642 : std_logic_vector(0 to 0) := (others => '0');
    variable r3641 : std_logic_vector(0 to 0) := (others => '0');
    variable r3640 : std_logic_vector(0 to 0) := (others => '0');
    variable r3639 : std_logic_vector(0 to 0) := (others => '0');
    variable r3638 : std_logic_vector(0 to 0) := (others => '0');
    variable r3637 : std_logic_vector(0 to 0) := (others => '0');
    variable r3636 : std_logic_vector(0 to 0) := (others => '0');
    variable r3635 : std_logic_vector(0 to 0) := (others => '0');
    variable r3634 : std_logic_vector(0 to 0) := (others => '0');
    variable r3633 : std_logic_vector(0 to 0) := (others => '0');
    variable r3632 : std_logic_vector(0 to 0) := (others => '0');
    variable r3631 : std_logic_vector(0 to 0) := (others => '0');
    variable r3630 : std_logic_vector(0 to 0) := (others => '0');
    variable r3629 : std_logic_vector(0 to 0) := (others => '0');
    variable r3628 : std_logic_vector(0 to 0) := (others => '0');
    variable r3627 : std_logic_vector(0 to 0) := (others => '0');
    variable r3626 : std_logic_vector(0 to 0) := (others => '0');
    variable r3625 : std_logic_vector(0 to 0) := (others => '0');
    variable r3624 : std_logic_vector(0 to 0) := (others => '0');
    variable r3623 : std_logic_vector(0 to 0) := (others => '0');
    variable r3622 : std_logic_vector(0 to 0) := (others => '0');
    variable r3621 : std_logic_vector(0 to 0) := (others => '0');
    variable r3620 : std_logic_vector(0 to 0) := (others => '0');
    variable r3619 : std_logic_vector(0 to 0) := (others => '0');
    variable r3618 : std_logic_vector(0 to 0) := (others => '0');
    variable r3617 : std_logic_vector(0 to 0) := (others => '0');
    variable r3616 : std_logic_vector(0 to 0) := (others => '0');
    variable r3615 : std_logic_vector(0 to 0) := (others => '0');
    variable r3614 : std_logic_vector(0 to 0) := (others => '0');
    variable r3613 : std_logic_vector(0 to 0) := (others => '0');
    variable r3612 : std_logic_vector(0 to 0) := (others => '0');
    variable r3611 : std_logic_vector(0 to 0) := (others => '0');
    variable r3610 : std_logic_vector(0 to 0) := (others => '0');
    variable r3609 : std_logic_vector(0 to 0) := (others => '0');
    variable r3608 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r3609 := "1";
    null;
    r3610 := (r3609);
    r3611 := "1";
    null;
    r3612 := (r3611);
    r3613 := "0";
    null;
    r3614 := (r3613);
    r3615 := "0";
    null;
    r3616 := (r3615);
    r3617 := "0";
    null;
    r3618 := (r3617);
    r3619 := "1";
    null;
    r3620 := (r3619);
    r3621 := "1";
    null;
    r3622 := (r3621);
    r3623 := "0";
    null;
    r3624 := (r3623);
    r3625 := "1";
    null;
    r3626 := (r3625);
    r3627 := "1";
    null;
    r3628 := (r3627);
    r3629 := "1";
    null;
    r3630 := (r3629);
    r3631 := "0";
    null;
    r3632 := (r3631);
    r3633 := "0";
    null;
    r3634 := (r3633);
    r3635 := "0";
    null;
    r3636 := (r3635);
    r3637 := "0";
    null;
    r3638 := (r3637);
    r3639 := "0";
    null;
    r3640 := (r3639);
    r3641 := "0";
    null;
    r3642 := (r3641);
    r3643 := "0";
    null;
    r3644 := (r3643);
    r3645 := "0";
    null;
    r3646 := (r3645);
    r3647 := "0";
    null;
    r3648 := (r3647);
    r3649 := "1";
    null;
    r3650 := (r3649);
    r3651 := "0";
    null;
    r3652 := (r3651);
    r3653 := "1";
    null;
    r3654 := (r3653);
    r3655 := "1";
    null;
    r3656 := (r3655);
    r3657 := "1";
    null;
    r3658 := (r3657);
    r3659 := "1";
    null;
    r3660 := (r3659);
    r3661 := "1";
    null;
    r3662 := (r3661);
    r3663 := "1";
    null;
    r3664 := (r3663);
    r3665 := "0";
    null;
    r3666 := (r3665);
    r3667 := "0";
    null;
    r3668 := (r3667);
    r3669 := "1";
    null;
    r3670 := (r3669);
    r3671 := "1";
    null;
    r3672 := (r3671);
    r3608 := (r3610 & r3612 & r3614 & r3616 & r3618 & r3620 & r3622 & r3624 & r3626 & r3628 & r3630 & r3632 & r3634 & r3636 & r3638 & r3640 & r3642 & r3644 & r3646 & r3648 & r3650 & r3652 & r3654 & r3656 & r3658 & r3660 & r3662 & r3664 & r3666 & r3668 & r3670 & r3672);
    return r3608;
  end rewire_MetaprogrammingRW.wc6e00bf3_3607;
  function rewire_MetaprogrammingRW.wbf597fc7_3538 return std_logic_vector
  is
    variable r3603 : std_logic_vector(0 to 0) := (others => '0');
    variable r3602 : std_logic_vector(0 to 0) := (others => '0');
    variable r3601 : std_logic_vector(0 to 0) := (others => '0');
    variable r3600 : std_logic_vector(0 to 0) := (others => '0');
    variable r3599 : std_logic_vector(0 to 0) := (others => '0');
    variable r3598 : std_logic_vector(0 to 0) := (others => '0');
    variable r3597 : std_logic_vector(0 to 0) := (others => '0');
    variable r3596 : std_logic_vector(0 to 0) := (others => '0');
    variable r3595 : std_logic_vector(0 to 0) := (others => '0');
    variable r3594 : std_logic_vector(0 to 0) := (others => '0');
    variable r3593 : std_logic_vector(0 to 0) := (others => '0');
    variable r3592 : std_logic_vector(0 to 0) := (others => '0');
    variable r3591 : std_logic_vector(0 to 0) := (others => '0');
    variable r3590 : std_logic_vector(0 to 0) := (others => '0');
    variable r3589 : std_logic_vector(0 to 0) := (others => '0');
    variable r3588 : std_logic_vector(0 to 0) := (others => '0');
    variable r3587 : std_logic_vector(0 to 0) := (others => '0');
    variable r3586 : std_logic_vector(0 to 0) := (others => '0');
    variable r3585 : std_logic_vector(0 to 0) := (others => '0');
    variable r3584 : std_logic_vector(0 to 0) := (others => '0');
    variable r3583 : std_logic_vector(0 to 0) := (others => '0');
    variable r3582 : std_logic_vector(0 to 0) := (others => '0');
    variable r3581 : std_logic_vector(0 to 0) := (others => '0');
    variable r3580 : std_logic_vector(0 to 0) := (others => '0');
    variable r3579 : std_logic_vector(0 to 0) := (others => '0');
    variable r3578 : std_logic_vector(0 to 0) := (others => '0');
    variable r3577 : std_logic_vector(0 to 0) := (others => '0');
    variable r3576 : std_logic_vector(0 to 0) := (others => '0');
    variable r3575 : std_logic_vector(0 to 0) := (others => '0');
    variable r3574 : std_logic_vector(0 to 0) := (others => '0');
    variable r3573 : std_logic_vector(0 to 0) := (others => '0');
    variable r3572 : std_logic_vector(0 to 0) := (others => '0');
    variable r3571 : std_logic_vector(0 to 0) := (others => '0');
    variable r3570 : std_logic_vector(0 to 0) := (others => '0');
    variable r3569 : std_logic_vector(0 to 0) := (others => '0');
    variable r3568 : std_logic_vector(0 to 0) := (others => '0');
    variable r3567 : std_logic_vector(0 to 0) := (others => '0');
    variable r3566 : std_logic_vector(0 to 0) := (others => '0');
    variable r3565 : std_logic_vector(0 to 0) := (others => '0');
    variable r3564 : std_logic_vector(0 to 0) := (others => '0');
    variable r3563 : std_logic_vector(0 to 0) := (others => '0');
    variable r3562 : std_logic_vector(0 to 0) := (others => '0');
    variable r3561 : std_logic_vector(0 to 0) := (others => '0');
    variable r3560 : std_logic_vector(0 to 0) := (others => '0');
    variable r3559 : std_logic_vector(0 to 0) := (others => '0');
    variable r3558 : std_logic_vector(0 to 0) := (others => '0');
    variable r3557 : std_logic_vector(0 to 0) := (others => '0');
    variable r3556 : std_logic_vector(0 to 0) := (others => '0');
    variable r3555 : std_logic_vector(0 to 0) := (others => '0');
    variable r3554 : std_logic_vector(0 to 0) := (others => '0');
    variable r3553 : std_logic_vector(0 to 0) := (others => '0');
    variable r3552 : std_logic_vector(0 to 0) := (others => '0');
    variable r3551 : std_logic_vector(0 to 0) := (others => '0');
    variable r3550 : std_logic_vector(0 to 0) := (others => '0');
    variable r3549 : std_logic_vector(0 to 0) := (others => '0');
    variable r3548 : std_logic_vector(0 to 0) := (others => '0');
    variable r3547 : std_logic_vector(0 to 0) := (others => '0');
    variable r3546 : std_logic_vector(0 to 0) := (others => '0');
    variable r3545 : std_logic_vector(0 to 0) := (others => '0');
    variable r3544 : std_logic_vector(0 to 0) := (others => '0');
    variable r3543 : std_logic_vector(0 to 0) := (others => '0');
    variable r3542 : std_logic_vector(0 to 0) := (others => '0');
    variable r3541 : std_logic_vector(0 to 0) := (others => '0');
    variable r3540 : std_logic_vector(0 to 0) := (others => '0');
    variable r3539 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r3540 := "1";
    null;
    r3541 := (r3540);
    r3542 := "0";
    null;
    r3543 := (r3542);
    r3544 := "1";
    null;
    r3545 := (r3544);
    r3546 := "1";
    null;
    r3547 := (r3546);
    r3548 := "1";
    null;
    r3549 := (r3548);
    r3550 := "1";
    null;
    r3551 := (r3550);
    r3552 := "1";
    null;
    r3553 := (r3552);
    r3554 := "1";
    null;
    r3555 := (r3554);
    r3556 := "0";
    null;
    r3557 := (r3556);
    r3558 := "1";
    null;
    r3559 := (r3558);
    r3560 := "0";
    null;
    r3561 := (r3560);
    r3562 := "1";
    null;
    r3563 := (r3562);
    r3564 := "1";
    null;
    r3565 := (r3564);
    r3566 := "0";
    null;
    r3567 := (r3566);
    r3568 := "0";
    null;
    r3569 := (r3568);
    r3570 := "1";
    null;
    r3571 := (r3570);
    r3572 := "0";
    null;
    r3573 := (r3572);
    r3574 := "1";
    null;
    r3575 := (r3574);
    r3576 := "1";
    null;
    r3577 := (r3576);
    r3578 := "1";
    null;
    r3579 := (r3578);
    r3580 := "1";
    null;
    r3581 := (r3580);
    r3582 := "1";
    null;
    r3583 := (r3582);
    r3584 := "1";
    null;
    r3585 := (r3584);
    r3586 := "1";
    null;
    r3587 := (r3586);
    r3588 := "1";
    null;
    r3589 := (r3588);
    r3590 := "1";
    null;
    r3591 := (r3590);
    r3592 := "0";
    null;
    r3593 := (r3592);
    r3594 := "0";
    null;
    r3595 := (r3594);
    r3596 := "0";
    null;
    r3597 := (r3596);
    r3598 := "1";
    null;
    r3599 := (r3598);
    r3600 := "1";
    null;
    r3601 := (r3600);
    r3602 := "1";
    null;
    r3603 := (r3602);
    r3539 := (r3541 & r3543 & r3545 & r3547 & r3549 & r3551 & r3553 & r3555 & r3557 & r3559 & r3561 & r3563 & r3565 & r3567 & r3569 & r3571 & r3573 & r3575 & r3577 & r3579 & r3581 & r3583 & r3585 & r3587 & r3589 & r3591 & r3593 & r3595 & r3597 & r3599 & r3601 & r3603);
    return r3539;
  end rewire_MetaprogrammingRW.wbf597fc7_3538;
  function rewire_MetaprogrammingRW.wb00327c8_3469 return std_logic_vector
  is
    variable r3534 : std_logic_vector(0 to 0) := (others => '0');
    variable r3533 : std_logic_vector(0 to 0) := (others => '0');
    variable r3532 : std_logic_vector(0 to 0) := (others => '0');
    variable r3531 : std_logic_vector(0 to 0) := (others => '0');
    variable r3530 : std_logic_vector(0 to 0) := (others => '0');
    variable r3529 : std_logic_vector(0 to 0) := (others => '0');
    variable r3528 : std_logic_vector(0 to 0) := (others => '0');
    variable r3527 : std_logic_vector(0 to 0) := (others => '0');
    variable r3526 : std_logic_vector(0 to 0) := (others => '0');
    variable r3525 : std_logic_vector(0 to 0) := (others => '0');
    variable r3524 : std_logic_vector(0 to 0) := (others => '0');
    variable r3523 : std_logic_vector(0 to 0) := (others => '0');
    variable r3522 : std_logic_vector(0 to 0) := (others => '0');
    variable r3521 : std_logic_vector(0 to 0) := (others => '0');
    variable r3520 : std_logic_vector(0 to 0) := (others => '0');
    variable r3519 : std_logic_vector(0 to 0) := (others => '0');
    variable r3518 : std_logic_vector(0 to 0) := (others => '0');
    variable r3517 : std_logic_vector(0 to 0) := (others => '0');
    variable r3516 : std_logic_vector(0 to 0) := (others => '0');
    variable r3515 : std_logic_vector(0 to 0) := (others => '0');
    variable r3514 : std_logic_vector(0 to 0) := (others => '0');
    variable r3513 : std_logic_vector(0 to 0) := (others => '0');
    variable r3512 : std_logic_vector(0 to 0) := (others => '0');
    variable r3511 : std_logic_vector(0 to 0) := (others => '0');
    variable r3510 : std_logic_vector(0 to 0) := (others => '0');
    variable r3509 : std_logic_vector(0 to 0) := (others => '0');
    variable r3508 : std_logic_vector(0 to 0) := (others => '0');
    variable r3507 : std_logic_vector(0 to 0) := (others => '0');
    variable r3506 : std_logic_vector(0 to 0) := (others => '0');
    variable r3505 : std_logic_vector(0 to 0) := (others => '0');
    variable r3504 : std_logic_vector(0 to 0) := (others => '0');
    variable r3503 : std_logic_vector(0 to 0) := (others => '0');
    variable r3502 : std_logic_vector(0 to 0) := (others => '0');
    variable r3501 : std_logic_vector(0 to 0) := (others => '0');
    variable r3500 : std_logic_vector(0 to 0) := (others => '0');
    variable r3499 : std_logic_vector(0 to 0) := (others => '0');
    variable r3498 : std_logic_vector(0 to 0) := (others => '0');
    variable r3497 : std_logic_vector(0 to 0) := (others => '0');
    variable r3496 : std_logic_vector(0 to 0) := (others => '0');
    variable r3495 : std_logic_vector(0 to 0) := (others => '0');
    variable r3494 : std_logic_vector(0 to 0) := (others => '0');
    variable r3493 : std_logic_vector(0 to 0) := (others => '0');
    variable r3492 : std_logic_vector(0 to 0) := (others => '0');
    variable r3491 : std_logic_vector(0 to 0) := (others => '0');
    variable r3490 : std_logic_vector(0 to 0) := (others => '0');
    variable r3489 : std_logic_vector(0 to 0) := (others => '0');
    variable r3488 : std_logic_vector(0 to 0) := (others => '0');
    variable r3487 : std_logic_vector(0 to 0) := (others => '0');
    variable r3486 : std_logic_vector(0 to 0) := (others => '0');
    variable r3485 : std_logic_vector(0 to 0) := (others => '0');
    variable r3484 : std_logic_vector(0 to 0) := (others => '0');
    variable r3483 : std_logic_vector(0 to 0) := (others => '0');
    variable r3482 : std_logic_vector(0 to 0) := (others => '0');
    variable r3481 : std_logic_vector(0 to 0) := (others => '0');
    variable r3480 : std_logic_vector(0 to 0) := (others => '0');
    variable r3479 : std_logic_vector(0 to 0) := (others => '0');
    variable r3478 : std_logic_vector(0 to 0) := (others => '0');
    variable r3477 : std_logic_vector(0 to 0) := (others => '0');
    variable r3476 : std_logic_vector(0 to 0) := (others => '0');
    variable r3475 : std_logic_vector(0 to 0) := (others => '0');
    variable r3474 : std_logic_vector(0 to 0) := (others => '0');
    variable r3473 : std_logic_vector(0 to 0) := (others => '0');
    variable r3472 : std_logic_vector(0 to 0) := (others => '0');
    variable r3471 : std_logic_vector(0 to 0) := (others => '0');
    variable r3470 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r3471 := "1";
    null;
    r3472 := (r3471);
    r3473 := "0";
    null;
    r3474 := (r3473);
    r3475 := "1";
    null;
    r3476 := (r3475);
    r3477 := "1";
    null;
    r3478 := (r3477);
    r3479 := "0";
    null;
    r3480 := (r3479);
    r3481 := "0";
    null;
    r3482 := (r3481);
    r3483 := "0";
    null;
    r3484 := (r3483);
    r3485 := "0";
    null;
    r3486 := (r3485);
    r3487 := "0";
    null;
    r3488 := (r3487);
    r3489 := "0";
    null;
    r3490 := (r3489);
    r3491 := "0";
    null;
    r3492 := (r3491);
    r3493 := "0";
    null;
    r3494 := (r3493);
    r3495 := "0";
    null;
    r3496 := (r3495);
    r3497 := "0";
    null;
    r3498 := (r3497);
    r3499 := "1";
    null;
    r3500 := (r3499);
    r3501 := "1";
    null;
    r3502 := (r3501);
    r3503 := "0";
    null;
    r3504 := (r3503);
    r3505 := "0";
    null;
    r3506 := (r3505);
    r3507 := "1";
    null;
    r3508 := (r3507);
    r3509 := "0";
    null;
    r3510 := (r3509);
    r3511 := "0";
    null;
    r3512 := (r3511);
    r3513 := "1";
    null;
    r3514 := (r3513);
    r3515 := "1";
    null;
    r3516 := (r3515);
    r3517 := "1";
    null;
    r3518 := (r3517);
    r3519 := "1";
    null;
    r3520 := (r3519);
    r3521 := "1";
    null;
    r3522 := (r3521);
    r3523 := "0";
    null;
    r3524 := (r3523);
    r3525 := "0";
    null;
    r3526 := (r3525);
    r3527 := "1";
    null;
    r3528 := (r3527);
    r3529 := "0";
    null;
    r3530 := (r3529);
    r3531 := "0";
    null;
    r3532 := (r3531);
    r3533 := "0";
    null;
    r3534 := (r3533);
    r3470 := (r3472 & r3474 & r3476 & r3478 & r3480 & r3482 & r3484 & r3486 & r3488 & r3490 & r3492 & r3494 & r3496 & r3498 & r3500 & r3502 & r3504 & r3506 & r3508 & r3510 & r3512 & r3514 & r3516 & r3518 & r3520 & r3522 & r3524 & r3526 & r3528 & r3530 & r3532 & r3534);
    return r3470;
  end rewire_MetaprogrammingRW.wb00327c8_3469;
  function rewire_MetaprogrammingRW.wa831c66d_3400 return std_logic_vector
  is
    variable r3465 : std_logic_vector(0 to 0) := (others => '0');
    variable r3464 : std_logic_vector(0 to 0) := (others => '0');
    variable r3463 : std_logic_vector(0 to 0) := (others => '0');
    variable r3462 : std_logic_vector(0 to 0) := (others => '0');
    variable r3461 : std_logic_vector(0 to 0) := (others => '0');
    variable r3460 : std_logic_vector(0 to 0) := (others => '0');
    variable r3459 : std_logic_vector(0 to 0) := (others => '0');
    variable r3458 : std_logic_vector(0 to 0) := (others => '0');
    variable r3457 : std_logic_vector(0 to 0) := (others => '0');
    variable r3456 : std_logic_vector(0 to 0) := (others => '0');
    variable r3455 : std_logic_vector(0 to 0) := (others => '0');
    variable r3454 : std_logic_vector(0 to 0) := (others => '0');
    variable r3453 : std_logic_vector(0 to 0) := (others => '0');
    variable r3452 : std_logic_vector(0 to 0) := (others => '0');
    variable r3451 : std_logic_vector(0 to 0) := (others => '0');
    variable r3450 : std_logic_vector(0 to 0) := (others => '0');
    variable r3449 : std_logic_vector(0 to 0) := (others => '0');
    variable r3448 : std_logic_vector(0 to 0) := (others => '0');
    variable r3447 : std_logic_vector(0 to 0) := (others => '0');
    variable r3446 : std_logic_vector(0 to 0) := (others => '0');
    variable r3445 : std_logic_vector(0 to 0) := (others => '0');
    variable r3444 : std_logic_vector(0 to 0) := (others => '0');
    variable r3443 : std_logic_vector(0 to 0) := (others => '0');
    variable r3442 : std_logic_vector(0 to 0) := (others => '0');
    variable r3441 : std_logic_vector(0 to 0) := (others => '0');
    variable r3440 : std_logic_vector(0 to 0) := (others => '0');
    variable r3439 : std_logic_vector(0 to 0) := (others => '0');
    variable r3438 : std_logic_vector(0 to 0) := (others => '0');
    variable r3437 : std_logic_vector(0 to 0) := (others => '0');
    variable r3436 : std_logic_vector(0 to 0) := (others => '0');
    variable r3435 : std_logic_vector(0 to 0) := (others => '0');
    variable r3434 : std_logic_vector(0 to 0) := (others => '0');
    variable r3433 : std_logic_vector(0 to 0) := (others => '0');
    variable r3432 : std_logic_vector(0 to 0) := (others => '0');
    variable r3431 : std_logic_vector(0 to 0) := (others => '0');
    variable r3430 : std_logic_vector(0 to 0) := (others => '0');
    variable r3429 : std_logic_vector(0 to 0) := (others => '0');
    variable r3428 : std_logic_vector(0 to 0) := (others => '0');
    variable r3427 : std_logic_vector(0 to 0) := (others => '0');
    variable r3426 : std_logic_vector(0 to 0) := (others => '0');
    variable r3425 : std_logic_vector(0 to 0) := (others => '0');
    variable r3424 : std_logic_vector(0 to 0) := (others => '0');
    variable r3423 : std_logic_vector(0 to 0) := (others => '0');
    variable r3422 : std_logic_vector(0 to 0) := (others => '0');
    variable r3421 : std_logic_vector(0 to 0) := (others => '0');
    variable r3420 : std_logic_vector(0 to 0) := (others => '0');
    variable r3419 : std_logic_vector(0 to 0) := (others => '0');
    variable r3418 : std_logic_vector(0 to 0) := (others => '0');
    variable r3417 : std_logic_vector(0 to 0) := (others => '0');
    variable r3416 : std_logic_vector(0 to 0) := (others => '0');
    variable r3415 : std_logic_vector(0 to 0) := (others => '0');
    variable r3414 : std_logic_vector(0 to 0) := (others => '0');
    variable r3413 : std_logic_vector(0 to 0) := (others => '0');
    variable r3412 : std_logic_vector(0 to 0) := (others => '0');
    variable r3411 : std_logic_vector(0 to 0) := (others => '0');
    variable r3410 : std_logic_vector(0 to 0) := (others => '0');
    variable r3409 : std_logic_vector(0 to 0) := (others => '0');
    variable r3408 : std_logic_vector(0 to 0) := (others => '0');
    variable r3407 : std_logic_vector(0 to 0) := (others => '0');
    variable r3406 : std_logic_vector(0 to 0) := (others => '0');
    variable r3405 : std_logic_vector(0 to 0) := (others => '0');
    variable r3404 : std_logic_vector(0 to 0) := (others => '0');
    variable r3403 : std_logic_vector(0 to 0) := (others => '0');
    variable r3402 : std_logic_vector(0 to 0) := (others => '0');
    variable r3401 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r3402 := "1";
    null;
    r3403 := (r3402);
    r3404 := "0";
    null;
    r3405 := (r3404);
    r3406 := "1";
    null;
    r3407 := (r3406);
    r3408 := "0";
    null;
    r3409 := (r3408);
    r3410 := "1";
    null;
    r3411 := (r3410);
    r3412 := "0";
    null;
    r3413 := (r3412);
    r3414 := "0";
    null;
    r3415 := (r3414);
    r3416 := "0";
    null;
    r3417 := (r3416);
    r3418 := "0";
    null;
    r3419 := (r3418);
    r3420 := "0";
    null;
    r3421 := (r3420);
    r3422 := "1";
    null;
    r3423 := (r3422);
    r3424 := "1";
    null;
    r3425 := (r3424);
    r3426 := "0";
    null;
    r3427 := (r3426);
    r3428 := "0";
    null;
    r3429 := (r3428);
    r3430 := "0";
    null;
    r3431 := (r3430);
    r3432 := "1";
    null;
    r3433 := (r3432);
    r3434 := "1";
    null;
    r3435 := (r3434);
    r3436 := "1";
    null;
    r3437 := (r3436);
    r3438 := "0";
    null;
    r3439 := (r3438);
    r3440 := "0";
    null;
    r3441 := (r3440);
    r3442 := "0";
    null;
    r3443 := (r3442);
    r3444 := "1";
    null;
    r3445 := (r3444);
    r3446 := "1";
    null;
    r3447 := (r3446);
    r3448 := "0";
    null;
    r3449 := (r3448);
    r3450 := "0";
    null;
    r3451 := (r3450);
    r3452 := "1";
    null;
    r3453 := (r3452);
    r3454 := "1";
    null;
    r3455 := (r3454);
    r3456 := "0";
    null;
    r3457 := (r3456);
    r3458 := "1";
    null;
    r3459 := (r3458);
    r3460 := "1";
    null;
    r3461 := (r3460);
    r3462 := "0";
    null;
    r3463 := (r3462);
    r3464 := "1";
    null;
    r3465 := (r3464);
    r3401 := (r3403 & r3405 & r3407 & r3409 & r3411 & r3413 & r3415 & r3417 & r3419 & r3421 & r3423 & r3425 & r3427 & r3429 & r3431 & r3433 & r3435 & r3437 & r3439 & r3441 & r3443 & r3445 & r3447 & r3449 & r3451 & r3453 & r3455 & r3457 & r3459 & r3461 & r3463 & r3465);
    return r3401;
  end rewire_MetaprogrammingRW.wa831c66d_3400;
  function rewire_MetaprogrammingRW.w983e5152_3331 return std_logic_vector
  is
    variable r3396 : std_logic_vector(0 to 0) := (others => '0');
    variable r3395 : std_logic_vector(0 to 0) := (others => '0');
    variable r3394 : std_logic_vector(0 to 0) := (others => '0');
    variable r3393 : std_logic_vector(0 to 0) := (others => '0');
    variable r3392 : std_logic_vector(0 to 0) := (others => '0');
    variable r3391 : std_logic_vector(0 to 0) := (others => '0');
    variable r3390 : std_logic_vector(0 to 0) := (others => '0');
    variable r3389 : std_logic_vector(0 to 0) := (others => '0');
    variable r3388 : std_logic_vector(0 to 0) := (others => '0');
    variable r3387 : std_logic_vector(0 to 0) := (others => '0');
    variable r3386 : std_logic_vector(0 to 0) := (others => '0');
    variable r3385 : std_logic_vector(0 to 0) := (others => '0');
    variable r3384 : std_logic_vector(0 to 0) := (others => '0');
    variable r3383 : std_logic_vector(0 to 0) := (others => '0');
    variable r3382 : std_logic_vector(0 to 0) := (others => '0');
    variable r3381 : std_logic_vector(0 to 0) := (others => '0');
    variable r3380 : std_logic_vector(0 to 0) := (others => '0');
    variable r3379 : std_logic_vector(0 to 0) := (others => '0');
    variable r3378 : std_logic_vector(0 to 0) := (others => '0');
    variable r3377 : std_logic_vector(0 to 0) := (others => '0');
    variable r3376 : std_logic_vector(0 to 0) := (others => '0');
    variable r3375 : std_logic_vector(0 to 0) := (others => '0');
    variable r3374 : std_logic_vector(0 to 0) := (others => '0');
    variable r3373 : std_logic_vector(0 to 0) := (others => '0');
    variable r3372 : std_logic_vector(0 to 0) := (others => '0');
    variable r3371 : std_logic_vector(0 to 0) := (others => '0');
    variable r3370 : std_logic_vector(0 to 0) := (others => '0');
    variable r3369 : std_logic_vector(0 to 0) := (others => '0');
    variable r3368 : std_logic_vector(0 to 0) := (others => '0');
    variable r3367 : std_logic_vector(0 to 0) := (others => '0');
    variable r3366 : std_logic_vector(0 to 0) := (others => '0');
    variable r3365 : std_logic_vector(0 to 0) := (others => '0');
    variable r3364 : std_logic_vector(0 to 0) := (others => '0');
    variable r3363 : std_logic_vector(0 to 0) := (others => '0');
    variable r3362 : std_logic_vector(0 to 0) := (others => '0');
    variable r3361 : std_logic_vector(0 to 0) := (others => '0');
    variable r3360 : std_logic_vector(0 to 0) := (others => '0');
    variable r3359 : std_logic_vector(0 to 0) := (others => '0');
    variable r3358 : std_logic_vector(0 to 0) := (others => '0');
    variable r3357 : std_logic_vector(0 to 0) := (others => '0');
    variable r3356 : std_logic_vector(0 to 0) := (others => '0');
    variable r3355 : std_logic_vector(0 to 0) := (others => '0');
    variable r3354 : std_logic_vector(0 to 0) := (others => '0');
    variable r3353 : std_logic_vector(0 to 0) := (others => '0');
    variable r3352 : std_logic_vector(0 to 0) := (others => '0');
    variable r3351 : std_logic_vector(0 to 0) := (others => '0');
    variable r3350 : std_logic_vector(0 to 0) := (others => '0');
    variable r3349 : std_logic_vector(0 to 0) := (others => '0');
    variable r3348 : std_logic_vector(0 to 0) := (others => '0');
    variable r3347 : std_logic_vector(0 to 0) := (others => '0');
    variable r3346 : std_logic_vector(0 to 0) := (others => '0');
    variable r3345 : std_logic_vector(0 to 0) := (others => '0');
    variable r3344 : std_logic_vector(0 to 0) := (others => '0');
    variable r3343 : std_logic_vector(0 to 0) := (others => '0');
    variable r3342 : std_logic_vector(0 to 0) := (others => '0');
    variable r3341 : std_logic_vector(0 to 0) := (others => '0');
    variable r3340 : std_logic_vector(0 to 0) := (others => '0');
    variable r3339 : std_logic_vector(0 to 0) := (others => '0');
    variable r3338 : std_logic_vector(0 to 0) := (others => '0');
    variable r3337 : std_logic_vector(0 to 0) := (others => '0');
    variable r3336 : std_logic_vector(0 to 0) := (others => '0');
    variable r3335 : std_logic_vector(0 to 0) := (others => '0');
    variable r3334 : std_logic_vector(0 to 0) := (others => '0');
    variable r3333 : std_logic_vector(0 to 0) := (others => '0');
    variable r3332 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r3333 := "1";
    null;
    r3334 := (r3333);
    r3335 := "0";
    null;
    r3336 := (r3335);
    r3337 := "0";
    null;
    r3338 := (r3337);
    r3339 := "1";
    null;
    r3340 := (r3339);
    r3341 := "1";
    null;
    r3342 := (r3341);
    r3343 := "0";
    null;
    r3344 := (r3343);
    r3345 := "0";
    null;
    r3346 := (r3345);
    r3347 := "0";
    null;
    r3348 := (r3347);
    r3349 := "0";
    null;
    r3350 := (r3349);
    r3351 := "0";
    null;
    r3352 := (r3351);
    r3353 := "1";
    null;
    r3354 := (r3353);
    r3355 := "1";
    null;
    r3356 := (r3355);
    r3357 := "1";
    null;
    r3358 := (r3357);
    r3359 := "1";
    null;
    r3360 := (r3359);
    r3361 := "1";
    null;
    r3362 := (r3361);
    r3363 := "0";
    null;
    r3364 := (r3363);
    r3365 := "0";
    null;
    r3366 := (r3365);
    r3367 := "1";
    null;
    r3368 := (r3367);
    r3369 := "0";
    null;
    r3370 := (r3369);
    r3371 := "1";
    null;
    r3372 := (r3371);
    r3373 := "0";
    null;
    r3374 := (r3373);
    r3375 := "0";
    null;
    r3376 := (r3375);
    r3377 := "0";
    null;
    r3378 := (r3377);
    r3379 := "1";
    null;
    r3380 := (r3379);
    r3381 := "0";
    null;
    r3382 := (r3381);
    r3383 := "1";
    null;
    r3384 := (r3383);
    r3385 := "0";
    null;
    r3386 := (r3385);
    r3387 := "1";
    null;
    r3388 := (r3387);
    r3389 := "0";
    null;
    r3390 := (r3389);
    r3391 := "0";
    null;
    r3392 := (r3391);
    r3393 := "1";
    null;
    r3394 := (r3393);
    r3395 := "0";
    null;
    r3396 := (r3395);
    r3332 := (r3334 & r3336 & r3338 & r3340 & r3342 & r3344 & r3346 & r3348 & r3350 & r3352 & r3354 & r3356 & r3358 & r3360 & r3362 & r3364 & r3366 & r3368 & r3370 & r3372 & r3374 & r3376 & r3378 & r3380 & r3382 & r3384 & r3386 & r3388 & r3390 & r3392 & r3394 & r3396);
    return r3332;
  end rewire_MetaprogrammingRW.w983e5152_3331;
  function rewire_MetaprogrammingRW.w76f988da_3262 return std_logic_vector
  is
    variable r3327 : std_logic_vector(0 to 0) := (others => '0');
    variable r3326 : std_logic_vector(0 to 0) := (others => '0');
    variable r3325 : std_logic_vector(0 to 0) := (others => '0');
    variable r3324 : std_logic_vector(0 to 0) := (others => '0');
    variable r3323 : std_logic_vector(0 to 0) := (others => '0');
    variable r3322 : std_logic_vector(0 to 0) := (others => '0');
    variable r3321 : std_logic_vector(0 to 0) := (others => '0');
    variable r3320 : std_logic_vector(0 to 0) := (others => '0');
    variable r3319 : std_logic_vector(0 to 0) := (others => '0');
    variable r3318 : std_logic_vector(0 to 0) := (others => '0');
    variable r3317 : std_logic_vector(0 to 0) := (others => '0');
    variable r3316 : std_logic_vector(0 to 0) := (others => '0');
    variable r3315 : std_logic_vector(0 to 0) := (others => '0');
    variable r3314 : std_logic_vector(0 to 0) := (others => '0');
    variable r3313 : std_logic_vector(0 to 0) := (others => '0');
    variable r3312 : std_logic_vector(0 to 0) := (others => '0');
    variable r3311 : std_logic_vector(0 to 0) := (others => '0');
    variable r3310 : std_logic_vector(0 to 0) := (others => '0');
    variable r3309 : std_logic_vector(0 to 0) := (others => '0');
    variable r3308 : std_logic_vector(0 to 0) := (others => '0');
    variable r3307 : std_logic_vector(0 to 0) := (others => '0');
    variable r3306 : std_logic_vector(0 to 0) := (others => '0');
    variable r3305 : std_logic_vector(0 to 0) := (others => '0');
    variable r3304 : std_logic_vector(0 to 0) := (others => '0');
    variable r3303 : std_logic_vector(0 to 0) := (others => '0');
    variable r3302 : std_logic_vector(0 to 0) := (others => '0');
    variable r3301 : std_logic_vector(0 to 0) := (others => '0');
    variable r3300 : std_logic_vector(0 to 0) := (others => '0');
    variable r3299 : std_logic_vector(0 to 0) := (others => '0');
    variable r3298 : std_logic_vector(0 to 0) := (others => '0');
    variable r3297 : std_logic_vector(0 to 0) := (others => '0');
    variable r3296 : std_logic_vector(0 to 0) := (others => '0');
    variable r3295 : std_logic_vector(0 to 0) := (others => '0');
    variable r3294 : std_logic_vector(0 to 0) := (others => '0');
    variable r3293 : std_logic_vector(0 to 0) := (others => '0');
    variable r3292 : std_logic_vector(0 to 0) := (others => '0');
    variable r3291 : std_logic_vector(0 to 0) := (others => '0');
    variable r3290 : std_logic_vector(0 to 0) := (others => '0');
    variable r3289 : std_logic_vector(0 to 0) := (others => '0');
    variable r3288 : std_logic_vector(0 to 0) := (others => '0');
    variable r3287 : std_logic_vector(0 to 0) := (others => '0');
    variable r3286 : std_logic_vector(0 to 0) := (others => '0');
    variable r3285 : std_logic_vector(0 to 0) := (others => '0');
    variable r3284 : std_logic_vector(0 to 0) := (others => '0');
    variable r3283 : std_logic_vector(0 to 0) := (others => '0');
    variable r3282 : std_logic_vector(0 to 0) := (others => '0');
    variable r3281 : std_logic_vector(0 to 0) := (others => '0');
    variable r3280 : std_logic_vector(0 to 0) := (others => '0');
    variable r3279 : std_logic_vector(0 to 0) := (others => '0');
    variable r3278 : std_logic_vector(0 to 0) := (others => '0');
    variable r3277 : std_logic_vector(0 to 0) := (others => '0');
    variable r3276 : std_logic_vector(0 to 0) := (others => '0');
    variable r3275 : std_logic_vector(0 to 0) := (others => '0');
    variable r3274 : std_logic_vector(0 to 0) := (others => '0');
    variable r3273 : std_logic_vector(0 to 0) := (others => '0');
    variable r3272 : std_logic_vector(0 to 0) := (others => '0');
    variable r3271 : std_logic_vector(0 to 0) := (others => '0');
    variable r3270 : std_logic_vector(0 to 0) := (others => '0');
    variable r3269 : std_logic_vector(0 to 0) := (others => '0');
    variable r3268 : std_logic_vector(0 to 0) := (others => '0');
    variable r3267 : std_logic_vector(0 to 0) := (others => '0');
    variable r3266 : std_logic_vector(0 to 0) := (others => '0');
    variable r3265 : std_logic_vector(0 to 0) := (others => '0');
    variable r3264 : std_logic_vector(0 to 0) := (others => '0');
    variable r3263 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r3264 := "0";
    null;
    r3265 := (r3264);
    r3266 := "1";
    null;
    r3267 := (r3266);
    r3268 := "1";
    null;
    r3269 := (r3268);
    r3270 := "1";
    null;
    r3271 := (r3270);
    r3272 := "0";
    null;
    r3273 := (r3272);
    r3274 := "1";
    null;
    r3275 := (r3274);
    r3276 := "1";
    null;
    r3277 := (r3276);
    r3278 := "0";
    null;
    r3279 := (r3278);
    r3280 := "1";
    null;
    r3281 := (r3280);
    r3282 := "1";
    null;
    r3283 := (r3282);
    r3284 := "1";
    null;
    r3285 := (r3284);
    r3286 := "1";
    null;
    r3287 := (r3286);
    r3288 := "1";
    null;
    r3289 := (r3288);
    r3290 := "0";
    null;
    r3291 := (r3290);
    r3292 := "0";
    null;
    r3293 := (r3292);
    r3294 := "1";
    null;
    r3295 := (r3294);
    r3296 := "1";
    null;
    r3297 := (r3296);
    r3298 := "0";
    null;
    r3299 := (r3298);
    r3300 := "0";
    null;
    r3301 := (r3300);
    r3302 := "0";
    null;
    r3303 := (r3302);
    r3304 := "1";
    null;
    r3305 := (r3304);
    r3306 := "0";
    null;
    r3307 := (r3306);
    r3308 := "0";
    null;
    r3309 := (r3308);
    r3310 := "0";
    null;
    r3311 := (r3310);
    r3312 := "1";
    null;
    r3313 := (r3312);
    r3314 := "1";
    null;
    r3315 := (r3314);
    r3316 := "0";
    null;
    r3317 := (r3316);
    r3318 := "1";
    null;
    r3319 := (r3318);
    r3320 := "1";
    null;
    r3321 := (r3320);
    r3322 := "0";
    null;
    r3323 := (r3322);
    r3324 := "1";
    null;
    r3325 := (r3324);
    r3326 := "0";
    null;
    r3327 := (r3326);
    r3263 := (r3265 & r3267 & r3269 & r3271 & r3273 & r3275 & r3277 & r3279 & r3281 & r3283 & r3285 & r3287 & r3289 & r3291 & r3293 & r3295 & r3297 & r3299 & r3301 & r3303 & r3305 & r3307 & r3309 & r3311 & r3313 & r3315 & r3317 & r3319 & r3321 & r3323 & r3325 & r3327);
    return r3263;
  end rewire_MetaprogrammingRW.w76f988da_3262;
  function rewire_MetaprogrammingRW.w5cb0a9dc_3193 return std_logic_vector
  is
    variable r3258 : std_logic_vector(0 to 0) := (others => '0');
    variable r3257 : std_logic_vector(0 to 0) := (others => '0');
    variable r3256 : std_logic_vector(0 to 0) := (others => '0');
    variable r3255 : std_logic_vector(0 to 0) := (others => '0');
    variable r3254 : std_logic_vector(0 to 0) := (others => '0');
    variable r3253 : std_logic_vector(0 to 0) := (others => '0');
    variable r3252 : std_logic_vector(0 to 0) := (others => '0');
    variable r3251 : std_logic_vector(0 to 0) := (others => '0');
    variable r3250 : std_logic_vector(0 to 0) := (others => '0');
    variable r3249 : std_logic_vector(0 to 0) := (others => '0');
    variable r3248 : std_logic_vector(0 to 0) := (others => '0');
    variable r3247 : std_logic_vector(0 to 0) := (others => '0');
    variable r3246 : std_logic_vector(0 to 0) := (others => '0');
    variable r3245 : std_logic_vector(0 to 0) := (others => '0');
    variable r3244 : std_logic_vector(0 to 0) := (others => '0');
    variable r3243 : std_logic_vector(0 to 0) := (others => '0');
    variable r3242 : std_logic_vector(0 to 0) := (others => '0');
    variable r3241 : std_logic_vector(0 to 0) := (others => '0');
    variable r3240 : std_logic_vector(0 to 0) := (others => '0');
    variable r3239 : std_logic_vector(0 to 0) := (others => '0');
    variable r3238 : std_logic_vector(0 to 0) := (others => '0');
    variable r3237 : std_logic_vector(0 to 0) := (others => '0');
    variable r3236 : std_logic_vector(0 to 0) := (others => '0');
    variable r3235 : std_logic_vector(0 to 0) := (others => '0');
    variable r3234 : std_logic_vector(0 to 0) := (others => '0');
    variable r3233 : std_logic_vector(0 to 0) := (others => '0');
    variable r3232 : std_logic_vector(0 to 0) := (others => '0');
    variable r3231 : std_logic_vector(0 to 0) := (others => '0');
    variable r3230 : std_logic_vector(0 to 0) := (others => '0');
    variable r3229 : std_logic_vector(0 to 0) := (others => '0');
    variable r3228 : std_logic_vector(0 to 0) := (others => '0');
    variable r3227 : std_logic_vector(0 to 0) := (others => '0');
    variable r3226 : std_logic_vector(0 to 0) := (others => '0');
    variable r3225 : std_logic_vector(0 to 0) := (others => '0');
    variable r3224 : std_logic_vector(0 to 0) := (others => '0');
    variable r3223 : std_logic_vector(0 to 0) := (others => '0');
    variable r3222 : std_logic_vector(0 to 0) := (others => '0');
    variable r3221 : std_logic_vector(0 to 0) := (others => '0');
    variable r3220 : std_logic_vector(0 to 0) := (others => '0');
    variable r3219 : std_logic_vector(0 to 0) := (others => '0');
    variable r3218 : std_logic_vector(0 to 0) := (others => '0');
    variable r3217 : std_logic_vector(0 to 0) := (others => '0');
    variable r3216 : std_logic_vector(0 to 0) := (others => '0');
    variable r3215 : std_logic_vector(0 to 0) := (others => '0');
    variable r3214 : std_logic_vector(0 to 0) := (others => '0');
    variable r3213 : std_logic_vector(0 to 0) := (others => '0');
    variable r3212 : std_logic_vector(0 to 0) := (others => '0');
    variable r3211 : std_logic_vector(0 to 0) := (others => '0');
    variable r3210 : std_logic_vector(0 to 0) := (others => '0');
    variable r3209 : std_logic_vector(0 to 0) := (others => '0');
    variable r3208 : std_logic_vector(0 to 0) := (others => '0');
    variable r3207 : std_logic_vector(0 to 0) := (others => '0');
    variable r3206 : std_logic_vector(0 to 0) := (others => '0');
    variable r3205 : std_logic_vector(0 to 0) := (others => '0');
    variable r3204 : std_logic_vector(0 to 0) := (others => '0');
    variable r3203 : std_logic_vector(0 to 0) := (others => '0');
    variable r3202 : std_logic_vector(0 to 0) := (others => '0');
    variable r3201 : std_logic_vector(0 to 0) := (others => '0');
    variable r3200 : std_logic_vector(0 to 0) := (others => '0');
    variable r3199 : std_logic_vector(0 to 0) := (others => '0');
    variable r3198 : std_logic_vector(0 to 0) := (others => '0');
    variable r3197 : std_logic_vector(0 to 0) := (others => '0');
    variable r3196 : std_logic_vector(0 to 0) := (others => '0');
    variable r3195 : std_logic_vector(0 to 0) := (others => '0');
    variable r3194 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r3195 := "0";
    null;
    r3196 := (r3195);
    r3197 := "1";
    null;
    r3198 := (r3197);
    r3199 := "0";
    null;
    r3200 := (r3199);
    r3201 := "1";
    null;
    r3202 := (r3201);
    r3203 := "1";
    null;
    r3204 := (r3203);
    r3205 := "1";
    null;
    r3206 := (r3205);
    r3207 := "0";
    null;
    r3208 := (r3207);
    r3209 := "0";
    null;
    r3210 := (r3209);
    r3211 := "1";
    null;
    r3212 := (r3211);
    r3213 := "0";
    null;
    r3214 := (r3213);
    r3215 := "1";
    null;
    r3216 := (r3215);
    r3217 := "1";
    null;
    r3218 := (r3217);
    r3219 := "0";
    null;
    r3220 := (r3219);
    r3221 := "0";
    null;
    r3222 := (r3221);
    r3223 := "0";
    null;
    r3224 := (r3223);
    r3225 := "0";
    null;
    r3226 := (r3225);
    r3227 := "1";
    null;
    r3228 := (r3227);
    r3229 := "0";
    null;
    r3230 := (r3229);
    r3231 := "1";
    null;
    r3232 := (r3231);
    r3233 := "0";
    null;
    r3234 := (r3233);
    r3235 := "1";
    null;
    r3236 := (r3235);
    r3237 := "0";
    null;
    r3238 := (r3237);
    r3239 := "0";
    null;
    r3240 := (r3239);
    r3241 := "1";
    null;
    r3242 := (r3241);
    r3243 := "1";
    null;
    r3244 := (r3243);
    r3245 := "1";
    null;
    r3246 := (r3245);
    r3247 := "0";
    null;
    r3248 := (r3247);
    r3249 := "1";
    null;
    r3250 := (r3249);
    r3251 := "1";
    null;
    r3252 := (r3251);
    r3253 := "1";
    null;
    r3254 := (r3253);
    r3255 := "0";
    null;
    r3256 := (r3255);
    r3257 := "0";
    null;
    r3258 := (r3257);
    r3194 := (r3196 & r3198 & r3200 & r3202 & r3204 & r3206 & r3208 & r3210 & r3212 & r3214 & r3216 & r3218 & r3220 & r3222 & r3224 & r3226 & r3228 & r3230 & r3232 & r3234 & r3236 & r3238 & r3240 & r3242 & r3244 & r3246 & r3248 & r3250 & r3252 & r3254 & r3256 & r3258);
    return r3194;
  end rewire_MetaprogrammingRW.w5cb0a9dc_3193;
  function rewire_MetaprogrammingRW.w4a7484aa_3124 return std_logic_vector
  is
    variable r3189 : std_logic_vector(0 to 0) := (others => '0');
    variable r3188 : std_logic_vector(0 to 0) := (others => '0');
    variable r3187 : std_logic_vector(0 to 0) := (others => '0');
    variable r3186 : std_logic_vector(0 to 0) := (others => '0');
    variable r3185 : std_logic_vector(0 to 0) := (others => '0');
    variable r3184 : std_logic_vector(0 to 0) := (others => '0');
    variable r3183 : std_logic_vector(0 to 0) := (others => '0');
    variable r3182 : std_logic_vector(0 to 0) := (others => '0');
    variable r3181 : std_logic_vector(0 to 0) := (others => '0');
    variable r3180 : std_logic_vector(0 to 0) := (others => '0');
    variable r3179 : std_logic_vector(0 to 0) := (others => '0');
    variable r3178 : std_logic_vector(0 to 0) := (others => '0');
    variable r3177 : std_logic_vector(0 to 0) := (others => '0');
    variable r3176 : std_logic_vector(0 to 0) := (others => '0');
    variable r3175 : std_logic_vector(0 to 0) := (others => '0');
    variable r3174 : std_logic_vector(0 to 0) := (others => '0');
    variable r3173 : std_logic_vector(0 to 0) := (others => '0');
    variable r3172 : std_logic_vector(0 to 0) := (others => '0');
    variable r3171 : std_logic_vector(0 to 0) := (others => '0');
    variable r3170 : std_logic_vector(0 to 0) := (others => '0');
    variable r3169 : std_logic_vector(0 to 0) := (others => '0');
    variable r3168 : std_logic_vector(0 to 0) := (others => '0');
    variable r3167 : std_logic_vector(0 to 0) := (others => '0');
    variable r3166 : std_logic_vector(0 to 0) := (others => '0');
    variable r3165 : std_logic_vector(0 to 0) := (others => '0');
    variable r3164 : std_logic_vector(0 to 0) := (others => '0');
    variable r3163 : std_logic_vector(0 to 0) := (others => '0');
    variable r3162 : std_logic_vector(0 to 0) := (others => '0');
    variable r3161 : std_logic_vector(0 to 0) := (others => '0');
    variable r3160 : std_logic_vector(0 to 0) := (others => '0');
    variable r3159 : std_logic_vector(0 to 0) := (others => '0');
    variable r3158 : std_logic_vector(0 to 0) := (others => '0');
    variable r3157 : std_logic_vector(0 to 0) := (others => '0');
    variable r3156 : std_logic_vector(0 to 0) := (others => '0');
    variable r3155 : std_logic_vector(0 to 0) := (others => '0');
    variable r3154 : std_logic_vector(0 to 0) := (others => '0');
    variable r3153 : std_logic_vector(0 to 0) := (others => '0');
    variable r3152 : std_logic_vector(0 to 0) := (others => '0');
    variable r3151 : std_logic_vector(0 to 0) := (others => '0');
    variable r3150 : std_logic_vector(0 to 0) := (others => '0');
    variable r3149 : std_logic_vector(0 to 0) := (others => '0');
    variable r3148 : std_logic_vector(0 to 0) := (others => '0');
    variable r3147 : std_logic_vector(0 to 0) := (others => '0');
    variable r3146 : std_logic_vector(0 to 0) := (others => '0');
    variable r3145 : std_logic_vector(0 to 0) := (others => '0');
    variable r3144 : std_logic_vector(0 to 0) := (others => '0');
    variable r3143 : std_logic_vector(0 to 0) := (others => '0');
    variable r3142 : std_logic_vector(0 to 0) := (others => '0');
    variable r3141 : std_logic_vector(0 to 0) := (others => '0');
    variable r3140 : std_logic_vector(0 to 0) := (others => '0');
    variable r3139 : std_logic_vector(0 to 0) := (others => '0');
    variable r3138 : std_logic_vector(0 to 0) := (others => '0');
    variable r3137 : std_logic_vector(0 to 0) := (others => '0');
    variable r3136 : std_logic_vector(0 to 0) := (others => '0');
    variable r3135 : std_logic_vector(0 to 0) := (others => '0');
    variable r3134 : std_logic_vector(0 to 0) := (others => '0');
    variable r3133 : std_logic_vector(0 to 0) := (others => '0');
    variable r3132 : std_logic_vector(0 to 0) := (others => '0');
    variable r3131 : std_logic_vector(0 to 0) := (others => '0');
    variable r3130 : std_logic_vector(0 to 0) := (others => '0');
    variable r3129 : std_logic_vector(0 to 0) := (others => '0');
    variable r3128 : std_logic_vector(0 to 0) := (others => '0');
    variable r3127 : std_logic_vector(0 to 0) := (others => '0');
    variable r3126 : std_logic_vector(0 to 0) := (others => '0');
    variable r3125 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r3126 := "0";
    null;
    r3127 := (r3126);
    r3128 := "1";
    null;
    r3129 := (r3128);
    r3130 := "0";
    null;
    r3131 := (r3130);
    r3132 := "0";
    null;
    r3133 := (r3132);
    r3134 := "1";
    null;
    r3135 := (r3134);
    r3136 := "0";
    null;
    r3137 := (r3136);
    r3138 := "1";
    null;
    r3139 := (r3138);
    r3140 := "0";
    null;
    r3141 := (r3140);
    r3142 := "0";
    null;
    r3143 := (r3142);
    r3144 := "1";
    null;
    r3145 := (r3144);
    r3146 := "1";
    null;
    r3147 := (r3146);
    r3148 := "1";
    null;
    r3149 := (r3148);
    r3150 := "0";
    null;
    r3151 := (r3150);
    r3152 := "1";
    null;
    r3153 := (r3152);
    r3154 := "0";
    null;
    r3155 := (r3154);
    r3156 := "0";
    null;
    r3157 := (r3156);
    r3158 := "1";
    null;
    r3159 := (r3158);
    r3160 := "0";
    null;
    r3161 := (r3160);
    r3162 := "0";
    null;
    r3163 := (r3162);
    r3164 := "0";
    null;
    r3165 := (r3164);
    r3166 := "0";
    null;
    r3167 := (r3166);
    r3168 := "1";
    null;
    r3169 := (r3168);
    r3170 := "0";
    null;
    r3171 := (r3170);
    r3172 := "0";
    null;
    r3173 := (r3172);
    r3174 := "1";
    null;
    r3175 := (r3174);
    r3176 := "0";
    null;
    r3177 := (r3176);
    r3178 := "1";
    null;
    r3179 := (r3178);
    r3180 := "0";
    null;
    r3181 := (r3180);
    r3182 := "1";
    null;
    r3183 := (r3182);
    r3184 := "0";
    null;
    r3185 := (r3184);
    r3186 := "1";
    null;
    r3187 := (r3186);
    r3188 := "0";
    null;
    r3189 := (r3188);
    r3125 := (r3127 & r3129 & r3131 & r3133 & r3135 & r3137 & r3139 & r3141 & r3143 & r3145 & r3147 & r3149 & r3151 & r3153 & r3155 & r3157 & r3159 & r3161 & r3163 & r3165 & r3167 & r3169 & r3171 & r3173 & r3175 & r3177 & r3179 & r3181 & r3183 & r3185 & r3187 & r3189);
    return r3125;
  end rewire_MetaprogrammingRW.w4a7484aa_3124;
  function rewire_MetaprogrammingRW.w2de92c6f_3055 return std_logic_vector
  is
    variable r3120 : std_logic_vector(0 to 0) := (others => '0');
    variable r3119 : std_logic_vector(0 to 0) := (others => '0');
    variable r3118 : std_logic_vector(0 to 0) := (others => '0');
    variable r3117 : std_logic_vector(0 to 0) := (others => '0');
    variable r3116 : std_logic_vector(0 to 0) := (others => '0');
    variable r3115 : std_logic_vector(0 to 0) := (others => '0');
    variable r3114 : std_logic_vector(0 to 0) := (others => '0');
    variable r3113 : std_logic_vector(0 to 0) := (others => '0');
    variable r3112 : std_logic_vector(0 to 0) := (others => '0');
    variable r3111 : std_logic_vector(0 to 0) := (others => '0');
    variable r3110 : std_logic_vector(0 to 0) := (others => '0');
    variable r3109 : std_logic_vector(0 to 0) := (others => '0');
    variable r3108 : std_logic_vector(0 to 0) := (others => '0');
    variable r3107 : std_logic_vector(0 to 0) := (others => '0');
    variable r3106 : std_logic_vector(0 to 0) := (others => '0');
    variable r3105 : std_logic_vector(0 to 0) := (others => '0');
    variable r3104 : std_logic_vector(0 to 0) := (others => '0');
    variable r3103 : std_logic_vector(0 to 0) := (others => '0');
    variable r3102 : std_logic_vector(0 to 0) := (others => '0');
    variable r3101 : std_logic_vector(0 to 0) := (others => '0');
    variable r3100 : std_logic_vector(0 to 0) := (others => '0');
    variable r3099 : std_logic_vector(0 to 0) := (others => '0');
    variable r3098 : std_logic_vector(0 to 0) := (others => '0');
    variable r3097 : std_logic_vector(0 to 0) := (others => '0');
    variable r3096 : std_logic_vector(0 to 0) := (others => '0');
    variable r3095 : std_logic_vector(0 to 0) := (others => '0');
    variable r3094 : std_logic_vector(0 to 0) := (others => '0');
    variable r3093 : std_logic_vector(0 to 0) := (others => '0');
    variable r3092 : std_logic_vector(0 to 0) := (others => '0');
    variable r3091 : std_logic_vector(0 to 0) := (others => '0');
    variable r3090 : std_logic_vector(0 to 0) := (others => '0');
    variable r3089 : std_logic_vector(0 to 0) := (others => '0');
    variable r3088 : std_logic_vector(0 to 0) := (others => '0');
    variable r3087 : std_logic_vector(0 to 0) := (others => '0');
    variable r3086 : std_logic_vector(0 to 0) := (others => '0');
    variable r3085 : std_logic_vector(0 to 0) := (others => '0');
    variable r3084 : std_logic_vector(0 to 0) := (others => '0');
    variable r3083 : std_logic_vector(0 to 0) := (others => '0');
    variable r3082 : std_logic_vector(0 to 0) := (others => '0');
    variable r3081 : std_logic_vector(0 to 0) := (others => '0');
    variable r3080 : std_logic_vector(0 to 0) := (others => '0');
    variable r3079 : std_logic_vector(0 to 0) := (others => '0');
    variable r3078 : std_logic_vector(0 to 0) := (others => '0');
    variable r3077 : std_logic_vector(0 to 0) := (others => '0');
    variable r3076 : std_logic_vector(0 to 0) := (others => '0');
    variable r3075 : std_logic_vector(0 to 0) := (others => '0');
    variable r3074 : std_logic_vector(0 to 0) := (others => '0');
    variable r3073 : std_logic_vector(0 to 0) := (others => '0');
    variable r3072 : std_logic_vector(0 to 0) := (others => '0');
    variable r3071 : std_logic_vector(0 to 0) := (others => '0');
    variable r3070 : std_logic_vector(0 to 0) := (others => '0');
    variable r3069 : std_logic_vector(0 to 0) := (others => '0');
    variable r3068 : std_logic_vector(0 to 0) := (others => '0');
    variable r3067 : std_logic_vector(0 to 0) := (others => '0');
    variable r3066 : std_logic_vector(0 to 0) := (others => '0');
    variable r3065 : std_logic_vector(0 to 0) := (others => '0');
    variable r3064 : std_logic_vector(0 to 0) := (others => '0');
    variable r3063 : std_logic_vector(0 to 0) := (others => '0');
    variable r3062 : std_logic_vector(0 to 0) := (others => '0');
    variable r3061 : std_logic_vector(0 to 0) := (others => '0');
    variable r3060 : std_logic_vector(0 to 0) := (others => '0');
    variable r3059 : std_logic_vector(0 to 0) := (others => '0');
    variable r3058 : std_logic_vector(0 to 0) := (others => '0');
    variable r3057 : std_logic_vector(0 to 0) := (others => '0');
    variable r3056 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r3057 := "0";
    null;
    r3058 := (r3057);
    r3059 := "0";
    null;
    r3060 := (r3059);
    r3061 := "1";
    null;
    r3062 := (r3061);
    r3063 := "0";
    null;
    r3064 := (r3063);
    r3065 := "1";
    null;
    r3066 := (r3065);
    r3067 := "1";
    null;
    r3068 := (r3067);
    r3069 := "0";
    null;
    r3070 := (r3069);
    r3071 := "1";
    null;
    r3072 := (r3071);
    r3073 := "1";
    null;
    r3074 := (r3073);
    r3075 := "1";
    null;
    r3076 := (r3075);
    r3077 := "1";
    null;
    r3078 := (r3077);
    r3079 := "0";
    null;
    r3080 := (r3079);
    r3081 := "1";
    null;
    r3082 := (r3081);
    r3083 := "0";
    null;
    r3084 := (r3083);
    r3085 := "0";
    null;
    r3086 := (r3085);
    r3087 := "1";
    null;
    r3088 := (r3087);
    r3089 := "0";
    null;
    r3090 := (r3089);
    r3091 := "0";
    null;
    r3092 := (r3091);
    r3093 := "1";
    null;
    r3094 := (r3093);
    r3095 := "0";
    null;
    r3096 := (r3095);
    r3097 := "1";
    null;
    r3098 := (r3097);
    r3099 := "1";
    null;
    r3100 := (r3099);
    r3101 := "0";
    null;
    r3102 := (r3101);
    r3103 := "0";
    null;
    r3104 := (r3103);
    r3105 := "0";
    null;
    r3106 := (r3105);
    r3107 := "1";
    null;
    r3108 := (r3107);
    r3109 := "1";
    null;
    r3110 := (r3109);
    r3111 := "0";
    null;
    r3112 := (r3111);
    r3113 := "1";
    null;
    r3114 := (r3113);
    r3115 := "1";
    null;
    r3116 := (r3115);
    r3117 := "1";
    null;
    r3118 := (r3117);
    r3119 := "1";
    null;
    r3120 := (r3119);
    r3056 := (r3058 & r3060 & r3062 & r3064 & r3066 & r3068 & r3070 & r3072 & r3074 & r3076 & r3078 & r3080 & r3082 & r3084 & r3086 & r3088 & r3090 & r3092 & r3094 & r3096 & r3098 & r3100 & r3102 & r3104 & r3106 & r3108 & r3110 & r3112 & r3114 & r3116 & r3118 & r3120);
    return r3056;
  end rewire_MetaprogrammingRW.w2de92c6f_3055;
  function rewire_MetaprogrammingRW.w240ca1cc_2986 return std_logic_vector
  is
    variable r3051 : std_logic_vector(0 to 0) := (others => '0');
    variable r3050 : std_logic_vector(0 to 0) := (others => '0');
    variable r3049 : std_logic_vector(0 to 0) := (others => '0');
    variable r3048 : std_logic_vector(0 to 0) := (others => '0');
    variable r3047 : std_logic_vector(0 to 0) := (others => '0');
    variable r3046 : std_logic_vector(0 to 0) := (others => '0');
    variable r3045 : std_logic_vector(0 to 0) := (others => '0');
    variable r3044 : std_logic_vector(0 to 0) := (others => '0');
    variable r3043 : std_logic_vector(0 to 0) := (others => '0');
    variable r3042 : std_logic_vector(0 to 0) := (others => '0');
    variable r3041 : std_logic_vector(0 to 0) := (others => '0');
    variable r3040 : std_logic_vector(0 to 0) := (others => '0');
    variable r3039 : std_logic_vector(0 to 0) := (others => '0');
    variable r3038 : std_logic_vector(0 to 0) := (others => '0');
    variable r3037 : std_logic_vector(0 to 0) := (others => '0');
    variable r3036 : std_logic_vector(0 to 0) := (others => '0');
    variable r3035 : std_logic_vector(0 to 0) := (others => '0');
    variable r3034 : std_logic_vector(0 to 0) := (others => '0');
    variable r3033 : std_logic_vector(0 to 0) := (others => '0');
    variable r3032 : std_logic_vector(0 to 0) := (others => '0');
    variable r3031 : std_logic_vector(0 to 0) := (others => '0');
    variable r3030 : std_logic_vector(0 to 0) := (others => '0');
    variable r3029 : std_logic_vector(0 to 0) := (others => '0');
    variable r3028 : std_logic_vector(0 to 0) := (others => '0');
    variable r3027 : std_logic_vector(0 to 0) := (others => '0');
    variable r3026 : std_logic_vector(0 to 0) := (others => '0');
    variable r3025 : std_logic_vector(0 to 0) := (others => '0');
    variable r3024 : std_logic_vector(0 to 0) := (others => '0');
    variable r3023 : std_logic_vector(0 to 0) := (others => '0');
    variable r3022 : std_logic_vector(0 to 0) := (others => '0');
    variable r3021 : std_logic_vector(0 to 0) := (others => '0');
    variable r3020 : std_logic_vector(0 to 0) := (others => '0');
    variable r3019 : std_logic_vector(0 to 0) := (others => '0');
    variable r3018 : std_logic_vector(0 to 0) := (others => '0');
    variable r3017 : std_logic_vector(0 to 0) := (others => '0');
    variable r3016 : std_logic_vector(0 to 0) := (others => '0');
    variable r3015 : std_logic_vector(0 to 0) := (others => '0');
    variable r3014 : std_logic_vector(0 to 0) := (others => '0');
    variable r3013 : std_logic_vector(0 to 0) := (others => '0');
    variable r3012 : std_logic_vector(0 to 0) := (others => '0');
    variable r3011 : std_logic_vector(0 to 0) := (others => '0');
    variable r3010 : std_logic_vector(0 to 0) := (others => '0');
    variable r3009 : std_logic_vector(0 to 0) := (others => '0');
    variable r3008 : std_logic_vector(0 to 0) := (others => '0');
    variable r3007 : std_logic_vector(0 to 0) := (others => '0');
    variable r3006 : std_logic_vector(0 to 0) := (others => '0');
    variable r3005 : std_logic_vector(0 to 0) := (others => '0');
    variable r3004 : std_logic_vector(0 to 0) := (others => '0');
    variable r3003 : std_logic_vector(0 to 0) := (others => '0');
    variable r3002 : std_logic_vector(0 to 0) := (others => '0');
    variable r3001 : std_logic_vector(0 to 0) := (others => '0');
    variable r3000 : std_logic_vector(0 to 0) := (others => '0');
    variable r2999 : std_logic_vector(0 to 0) := (others => '0');
    variable r2998 : std_logic_vector(0 to 0) := (others => '0');
    variable r2997 : std_logic_vector(0 to 0) := (others => '0');
    variable r2996 : std_logic_vector(0 to 0) := (others => '0');
    variable r2995 : std_logic_vector(0 to 0) := (others => '0');
    variable r2994 : std_logic_vector(0 to 0) := (others => '0');
    variable r2993 : std_logic_vector(0 to 0) := (others => '0');
    variable r2992 : std_logic_vector(0 to 0) := (others => '0');
    variable r2991 : std_logic_vector(0 to 0) := (others => '0');
    variable r2990 : std_logic_vector(0 to 0) := (others => '0');
    variable r2989 : std_logic_vector(0 to 0) := (others => '0');
    variable r2988 : std_logic_vector(0 to 0) := (others => '0');
    variable r2987 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r2988 := "0";
    null;
    r2989 := (r2988);
    r2990 := "0";
    null;
    r2991 := (r2990);
    r2992 := "1";
    null;
    r2993 := (r2992);
    r2994 := "0";
    null;
    r2995 := (r2994);
    r2996 := "0";
    null;
    r2997 := (r2996);
    r2998 := "1";
    null;
    r2999 := (r2998);
    r3000 := "0";
    null;
    r3001 := (r3000);
    r3002 := "0";
    null;
    r3003 := (r3002);
    r3004 := "0";
    null;
    r3005 := (r3004);
    r3006 := "0";
    null;
    r3007 := (r3006);
    r3008 := "0";
    null;
    r3009 := (r3008);
    r3010 := "0";
    null;
    r3011 := (r3010);
    r3012 := "1";
    null;
    r3013 := (r3012);
    r3014 := "1";
    null;
    r3015 := (r3014);
    r3016 := "0";
    null;
    r3017 := (r3016);
    r3018 := "0";
    null;
    r3019 := (r3018);
    r3020 := "1";
    null;
    r3021 := (r3020);
    r3022 := "0";
    null;
    r3023 := (r3022);
    r3024 := "1";
    null;
    r3025 := (r3024);
    r3026 := "0";
    null;
    r3027 := (r3026);
    r3028 := "0";
    null;
    r3029 := (r3028);
    r3030 := "0";
    null;
    r3031 := (r3030);
    r3032 := "0";
    null;
    r3033 := (r3032);
    r3034 := "1";
    null;
    r3035 := (r3034);
    r3036 := "1";
    null;
    r3037 := (r3036);
    r3038 := "1";
    null;
    r3039 := (r3038);
    r3040 := "0";
    null;
    r3041 := (r3040);
    r3042 := "0";
    null;
    r3043 := (r3042);
    r3044 := "1";
    null;
    r3045 := (r3044);
    r3046 := "1";
    null;
    r3047 := (r3046);
    r3048 := "0";
    null;
    r3049 := (r3048);
    r3050 := "0";
    null;
    r3051 := (r3050);
    r2987 := (r2989 & r2991 & r2993 & r2995 & r2997 & r2999 & r3001 & r3003 & r3005 & r3007 & r3009 & r3011 & r3013 & r3015 & r3017 & r3019 & r3021 & r3023 & r3025 & r3027 & r3029 & r3031 & r3033 & r3035 & r3037 & r3039 & r3041 & r3043 & r3045 & r3047 & r3049 & r3051);
    return r2987;
  end rewire_MetaprogrammingRW.w240ca1cc_2986;
  function rewire_MetaprogrammingRW.w0fc19dc6_2917 return std_logic_vector
  is
    variable r2982 : std_logic_vector(0 to 0) := (others => '0');
    variable r2981 : std_logic_vector(0 to 0) := (others => '0');
    variable r2980 : std_logic_vector(0 to 0) := (others => '0');
    variable r2979 : std_logic_vector(0 to 0) := (others => '0');
    variable r2978 : std_logic_vector(0 to 0) := (others => '0');
    variable r2977 : std_logic_vector(0 to 0) := (others => '0');
    variable r2976 : std_logic_vector(0 to 0) := (others => '0');
    variable r2975 : std_logic_vector(0 to 0) := (others => '0');
    variable r2974 : std_logic_vector(0 to 0) := (others => '0');
    variable r2973 : std_logic_vector(0 to 0) := (others => '0');
    variable r2972 : std_logic_vector(0 to 0) := (others => '0');
    variable r2971 : std_logic_vector(0 to 0) := (others => '0');
    variable r2970 : std_logic_vector(0 to 0) := (others => '0');
    variable r2969 : std_logic_vector(0 to 0) := (others => '0');
    variable r2968 : std_logic_vector(0 to 0) := (others => '0');
    variable r2967 : std_logic_vector(0 to 0) := (others => '0');
    variable r2966 : std_logic_vector(0 to 0) := (others => '0');
    variable r2965 : std_logic_vector(0 to 0) := (others => '0');
    variable r2964 : std_logic_vector(0 to 0) := (others => '0');
    variable r2963 : std_logic_vector(0 to 0) := (others => '0');
    variable r2962 : std_logic_vector(0 to 0) := (others => '0');
    variable r2961 : std_logic_vector(0 to 0) := (others => '0');
    variable r2960 : std_logic_vector(0 to 0) := (others => '0');
    variable r2959 : std_logic_vector(0 to 0) := (others => '0');
    variable r2958 : std_logic_vector(0 to 0) := (others => '0');
    variable r2957 : std_logic_vector(0 to 0) := (others => '0');
    variable r2956 : std_logic_vector(0 to 0) := (others => '0');
    variable r2955 : std_logic_vector(0 to 0) := (others => '0');
    variable r2954 : std_logic_vector(0 to 0) := (others => '0');
    variable r2953 : std_logic_vector(0 to 0) := (others => '0');
    variable r2952 : std_logic_vector(0 to 0) := (others => '0');
    variable r2951 : std_logic_vector(0 to 0) := (others => '0');
    variable r2950 : std_logic_vector(0 to 0) := (others => '0');
    variable r2949 : std_logic_vector(0 to 0) := (others => '0');
    variable r2948 : std_logic_vector(0 to 0) := (others => '0');
    variable r2947 : std_logic_vector(0 to 0) := (others => '0');
    variable r2946 : std_logic_vector(0 to 0) := (others => '0');
    variable r2945 : std_logic_vector(0 to 0) := (others => '0');
    variable r2944 : std_logic_vector(0 to 0) := (others => '0');
    variable r2943 : std_logic_vector(0 to 0) := (others => '0');
    variable r2942 : std_logic_vector(0 to 0) := (others => '0');
    variable r2941 : std_logic_vector(0 to 0) := (others => '0');
    variable r2940 : std_logic_vector(0 to 0) := (others => '0');
    variable r2939 : std_logic_vector(0 to 0) := (others => '0');
    variable r2938 : std_logic_vector(0 to 0) := (others => '0');
    variable r2937 : std_logic_vector(0 to 0) := (others => '0');
    variable r2936 : std_logic_vector(0 to 0) := (others => '0');
    variable r2935 : std_logic_vector(0 to 0) := (others => '0');
    variable r2934 : std_logic_vector(0 to 0) := (others => '0');
    variable r2933 : std_logic_vector(0 to 0) := (others => '0');
    variable r2932 : std_logic_vector(0 to 0) := (others => '0');
    variable r2931 : std_logic_vector(0 to 0) := (others => '0');
    variable r2930 : std_logic_vector(0 to 0) := (others => '0');
    variable r2929 : std_logic_vector(0 to 0) := (others => '0');
    variable r2928 : std_logic_vector(0 to 0) := (others => '0');
    variable r2927 : std_logic_vector(0 to 0) := (others => '0');
    variable r2926 : std_logic_vector(0 to 0) := (others => '0');
    variable r2925 : std_logic_vector(0 to 0) := (others => '0');
    variable r2924 : std_logic_vector(0 to 0) := (others => '0');
    variable r2923 : std_logic_vector(0 to 0) := (others => '0');
    variable r2922 : std_logic_vector(0 to 0) := (others => '0');
    variable r2921 : std_logic_vector(0 to 0) := (others => '0');
    variable r2920 : std_logic_vector(0 to 0) := (others => '0');
    variable r2919 : std_logic_vector(0 to 0) := (others => '0');
    variable r2918 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r2919 := "0";
    null;
    r2920 := (r2919);
    r2921 := "0";
    null;
    r2922 := (r2921);
    r2923 := "0";
    null;
    r2924 := (r2923);
    r2925 := "0";
    null;
    r2926 := (r2925);
    r2927 := "1";
    null;
    r2928 := (r2927);
    r2929 := "1";
    null;
    r2930 := (r2929);
    r2931 := "1";
    null;
    r2932 := (r2931);
    r2933 := "1";
    null;
    r2934 := (r2933);
    r2935 := "1";
    null;
    r2936 := (r2935);
    r2937 := "1";
    null;
    r2938 := (r2937);
    r2939 := "0";
    null;
    r2940 := (r2939);
    r2941 := "0";
    null;
    r2942 := (r2941);
    r2943 := "0";
    null;
    r2944 := (r2943);
    r2945 := "0";
    null;
    r2946 := (r2945);
    r2947 := "0";
    null;
    r2948 := (r2947);
    r2949 := "1";
    null;
    r2950 := (r2949);
    r2951 := "1";
    null;
    r2952 := (r2951);
    r2953 := "0";
    null;
    r2954 := (r2953);
    r2955 := "0";
    null;
    r2956 := (r2955);
    r2957 := "1";
    null;
    r2958 := (r2957);
    r2959 := "1";
    null;
    r2960 := (r2959);
    r2961 := "1";
    null;
    r2962 := (r2961);
    r2963 := "0";
    null;
    r2964 := (r2963);
    r2965 := "1";
    null;
    r2966 := (r2965);
    r2967 := "1";
    null;
    r2968 := (r2967);
    r2969 := "1";
    null;
    r2970 := (r2969);
    r2971 := "0";
    null;
    r2972 := (r2971);
    r2973 := "0";
    null;
    r2974 := (r2973);
    r2975 := "0";
    null;
    r2976 := (r2975);
    r2977 := "1";
    null;
    r2978 := (r2977);
    r2979 := "1";
    null;
    r2980 := (r2979);
    r2981 := "0";
    null;
    r2982 := (r2981);
    r2918 := (r2920 & r2922 & r2924 & r2926 & r2928 & r2930 & r2932 & r2934 & r2936 & r2938 & r2940 & r2942 & r2944 & r2946 & r2948 & r2950 & r2952 & r2954 & r2956 & r2958 & r2960 & r2962 & r2964 & r2966 & r2968 & r2970 & r2972 & r2974 & r2976 & r2978 & r2980 & r2982);
    return r2918;
  end rewire_MetaprogrammingRW.w0fc19dc6_2917;
  function rewire_MetaprogrammingRW.wefbe4786_2848 return std_logic_vector
  is
    variable r2913 : std_logic_vector(0 to 0) := (others => '0');
    variable r2912 : std_logic_vector(0 to 0) := (others => '0');
    variable r2911 : std_logic_vector(0 to 0) := (others => '0');
    variable r2910 : std_logic_vector(0 to 0) := (others => '0');
    variable r2909 : std_logic_vector(0 to 0) := (others => '0');
    variable r2908 : std_logic_vector(0 to 0) := (others => '0');
    variable r2907 : std_logic_vector(0 to 0) := (others => '0');
    variable r2906 : std_logic_vector(0 to 0) := (others => '0');
    variable r2905 : std_logic_vector(0 to 0) := (others => '0');
    variable r2904 : std_logic_vector(0 to 0) := (others => '0');
    variable r2903 : std_logic_vector(0 to 0) := (others => '0');
    variable r2902 : std_logic_vector(0 to 0) := (others => '0');
    variable r2901 : std_logic_vector(0 to 0) := (others => '0');
    variable r2900 : std_logic_vector(0 to 0) := (others => '0');
    variable r2899 : std_logic_vector(0 to 0) := (others => '0');
    variable r2898 : std_logic_vector(0 to 0) := (others => '0');
    variable r2897 : std_logic_vector(0 to 0) := (others => '0');
    variable r2896 : std_logic_vector(0 to 0) := (others => '0');
    variable r2895 : std_logic_vector(0 to 0) := (others => '0');
    variable r2894 : std_logic_vector(0 to 0) := (others => '0');
    variable r2893 : std_logic_vector(0 to 0) := (others => '0');
    variable r2892 : std_logic_vector(0 to 0) := (others => '0');
    variable r2891 : std_logic_vector(0 to 0) := (others => '0');
    variable r2890 : std_logic_vector(0 to 0) := (others => '0');
    variable r2889 : std_logic_vector(0 to 0) := (others => '0');
    variable r2888 : std_logic_vector(0 to 0) := (others => '0');
    variable r2887 : std_logic_vector(0 to 0) := (others => '0');
    variable r2886 : std_logic_vector(0 to 0) := (others => '0');
    variable r2885 : std_logic_vector(0 to 0) := (others => '0');
    variable r2884 : std_logic_vector(0 to 0) := (others => '0');
    variable r2883 : std_logic_vector(0 to 0) := (others => '0');
    variable r2882 : std_logic_vector(0 to 0) := (others => '0');
    variable r2881 : std_logic_vector(0 to 0) := (others => '0');
    variable r2880 : std_logic_vector(0 to 0) := (others => '0');
    variable r2879 : std_logic_vector(0 to 0) := (others => '0');
    variable r2878 : std_logic_vector(0 to 0) := (others => '0');
    variable r2877 : std_logic_vector(0 to 0) := (others => '0');
    variable r2876 : std_logic_vector(0 to 0) := (others => '0');
    variable r2875 : std_logic_vector(0 to 0) := (others => '0');
    variable r2874 : std_logic_vector(0 to 0) := (others => '0');
    variable r2873 : std_logic_vector(0 to 0) := (others => '0');
    variable r2872 : std_logic_vector(0 to 0) := (others => '0');
    variable r2871 : std_logic_vector(0 to 0) := (others => '0');
    variable r2870 : std_logic_vector(0 to 0) := (others => '0');
    variable r2869 : std_logic_vector(0 to 0) := (others => '0');
    variable r2868 : std_logic_vector(0 to 0) := (others => '0');
    variable r2867 : std_logic_vector(0 to 0) := (others => '0');
    variable r2866 : std_logic_vector(0 to 0) := (others => '0');
    variable r2865 : std_logic_vector(0 to 0) := (others => '0');
    variable r2864 : std_logic_vector(0 to 0) := (others => '0');
    variable r2863 : std_logic_vector(0 to 0) := (others => '0');
    variable r2862 : std_logic_vector(0 to 0) := (others => '0');
    variable r2861 : std_logic_vector(0 to 0) := (others => '0');
    variable r2860 : std_logic_vector(0 to 0) := (others => '0');
    variable r2859 : std_logic_vector(0 to 0) := (others => '0');
    variable r2858 : std_logic_vector(0 to 0) := (others => '0');
    variable r2857 : std_logic_vector(0 to 0) := (others => '0');
    variable r2856 : std_logic_vector(0 to 0) := (others => '0');
    variable r2855 : std_logic_vector(0 to 0) := (others => '0');
    variable r2854 : std_logic_vector(0 to 0) := (others => '0');
    variable r2853 : std_logic_vector(0 to 0) := (others => '0');
    variable r2852 : std_logic_vector(0 to 0) := (others => '0');
    variable r2851 : std_logic_vector(0 to 0) := (others => '0');
    variable r2850 : std_logic_vector(0 to 0) := (others => '0');
    variable r2849 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r2850 := "1";
    null;
    r2851 := (r2850);
    r2852 := "1";
    null;
    r2853 := (r2852);
    r2854 := "1";
    null;
    r2855 := (r2854);
    r2856 := "0";
    null;
    r2857 := (r2856);
    r2858 := "1";
    null;
    r2859 := (r2858);
    r2860 := "1";
    null;
    r2861 := (r2860);
    r2862 := "1";
    null;
    r2863 := (r2862);
    r2864 := "1";
    null;
    r2865 := (r2864);
    r2866 := "1";
    null;
    r2867 := (r2866);
    r2868 := "0";
    null;
    r2869 := (r2868);
    r2870 := "1";
    null;
    r2871 := (r2870);
    r2872 := "1";
    null;
    r2873 := (r2872);
    r2874 := "1";
    null;
    r2875 := (r2874);
    r2876 := "1";
    null;
    r2877 := (r2876);
    r2878 := "1";
    null;
    r2879 := (r2878);
    r2880 := "0";
    null;
    r2881 := (r2880);
    r2882 := "0";
    null;
    r2883 := (r2882);
    r2884 := "1";
    null;
    r2885 := (r2884);
    r2886 := "0";
    null;
    r2887 := (r2886);
    r2888 := "0";
    null;
    r2889 := (r2888);
    r2890 := "0";
    null;
    r2891 := (r2890);
    r2892 := "1";
    null;
    r2893 := (r2892);
    r2894 := "1";
    null;
    r2895 := (r2894);
    r2896 := "1";
    null;
    r2897 := (r2896);
    r2898 := "1";
    null;
    r2899 := (r2898);
    r2900 := "0";
    null;
    r2901 := (r2900);
    r2902 := "0";
    null;
    r2903 := (r2902);
    r2904 := "0";
    null;
    r2905 := (r2904);
    r2906 := "0";
    null;
    r2907 := (r2906);
    r2908 := "1";
    null;
    r2909 := (r2908);
    r2910 := "1";
    null;
    r2911 := (r2910);
    r2912 := "0";
    null;
    r2913 := (r2912);
    r2849 := (r2851 & r2853 & r2855 & r2857 & r2859 & r2861 & r2863 & r2865 & r2867 & r2869 & r2871 & r2873 & r2875 & r2877 & r2879 & r2881 & r2883 & r2885 & r2887 & r2889 & r2891 & r2893 & r2895 & r2897 & r2899 & r2901 & r2903 & r2905 & r2907 & r2909 & r2911 & r2913);
    return r2849;
  end rewire_MetaprogrammingRW.wefbe4786_2848;
  function rewire_MetaprogrammingRW.we49b69c1_2779 return std_logic_vector
  is
    variable r2844 : std_logic_vector(0 to 0) := (others => '0');
    variable r2843 : std_logic_vector(0 to 0) := (others => '0');
    variable r2842 : std_logic_vector(0 to 0) := (others => '0');
    variable r2841 : std_logic_vector(0 to 0) := (others => '0');
    variable r2840 : std_logic_vector(0 to 0) := (others => '0');
    variable r2839 : std_logic_vector(0 to 0) := (others => '0');
    variable r2838 : std_logic_vector(0 to 0) := (others => '0');
    variable r2837 : std_logic_vector(0 to 0) := (others => '0');
    variable r2836 : std_logic_vector(0 to 0) := (others => '0');
    variable r2835 : std_logic_vector(0 to 0) := (others => '0');
    variable r2834 : std_logic_vector(0 to 0) := (others => '0');
    variable r2833 : std_logic_vector(0 to 0) := (others => '0');
    variable r2832 : std_logic_vector(0 to 0) := (others => '0');
    variable r2831 : std_logic_vector(0 to 0) := (others => '0');
    variable r2830 : std_logic_vector(0 to 0) := (others => '0');
    variable r2829 : std_logic_vector(0 to 0) := (others => '0');
    variable r2828 : std_logic_vector(0 to 0) := (others => '0');
    variable r2827 : std_logic_vector(0 to 0) := (others => '0');
    variable r2826 : std_logic_vector(0 to 0) := (others => '0');
    variable r2825 : std_logic_vector(0 to 0) := (others => '0');
    variable r2824 : std_logic_vector(0 to 0) := (others => '0');
    variable r2823 : std_logic_vector(0 to 0) := (others => '0');
    variable r2822 : std_logic_vector(0 to 0) := (others => '0');
    variable r2821 : std_logic_vector(0 to 0) := (others => '0');
    variable r2820 : std_logic_vector(0 to 0) := (others => '0');
    variable r2819 : std_logic_vector(0 to 0) := (others => '0');
    variable r2818 : std_logic_vector(0 to 0) := (others => '0');
    variable r2817 : std_logic_vector(0 to 0) := (others => '0');
    variable r2816 : std_logic_vector(0 to 0) := (others => '0');
    variable r2815 : std_logic_vector(0 to 0) := (others => '0');
    variable r2814 : std_logic_vector(0 to 0) := (others => '0');
    variable r2813 : std_logic_vector(0 to 0) := (others => '0');
    variable r2812 : std_logic_vector(0 to 0) := (others => '0');
    variable r2811 : std_logic_vector(0 to 0) := (others => '0');
    variable r2810 : std_logic_vector(0 to 0) := (others => '0');
    variable r2809 : std_logic_vector(0 to 0) := (others => '0');
    variable r2808 : std_logic_vector(0 to 0) := (others => '0');
    variable r2807 : std_logic_vector(0 to 0) := (others => '0');
    variable r2806 : std_logic_vector(0 to 0) := (others => '0');
    variable r2805 : std_logic_vector(0 to 0) := (others => '0');
    variable r2804 : std_logic_vector(0 to 0) := (others => '0');
    variable r2803 : std_logic_vector(0 to 0) := (others => '0');
    variable r2802 : std_logic_vector(0 to 0) := (others => '0');
    variable r2801 : std_logic_vector(0 to 0) := (others => '0');
    variable r2800 : std_logic_vector(0 to 0) := (others => '0');
    variable r2799 : std_logic_vector(0 to 0) := (others => '0');
    variable r2798 : std_logic_vector(0 to 0) := (others => '0');
    variable r2797 : std_logic_vector(0 to 0) := (others => '0');
    variable r2796 : std_logic_vector(0 to 0) := (others => '0');
    variable r2795 : std_logic_vector(0 to 0) := (others => '0');
    variable r2794 : std_logic_vector(0 to 0) := (others => '0');
    variable r2793 : std_logic_vector(0 to 0) := (others => '0');
    variable r2792 : std_logic_vector(0 to 0) := (others => '0');
    variable r2791 : std_logic_vector(0 to 0) := (others => '0');
    variable r2790 : std_logic_vector(0 to 0) := (others => '0');
    variable r2789 : std_logic_vector(0 to 0) := (others => '0');
    variable r2788 : std_logic_vector(0 to 0) := (others => '0');
    variable r2787 : std_logic_vector(0 to 0) := (others => '0');
    variable r2786 : std_logic_vector(0 to 0) := (others => '0');
    variable r2785 : std_logic_vector(0 to 0) := (others => '0');
    variable r2784 : std_logic_vector(0 to 0) := (others => '0');
    variable r2783 : std_logic_vector(0 to 0) := (others => '0');
    variable r2782 : std_logic_vector(0 to 0) := (others => '0');
    variable r2781 : std_logic_vector(0 to 0) := (others => '0');
    variable r2780 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r2781 := "1";
    null;
    r2782 := (r2781);
    r2783 := "1";
    null;
    r2784 := (r2783);
    r2785 := "1";
    null;
    r2786 := (r2785);
    r2787 := "0";
    null;
    r2788 := (r2787);
    r2789 := "0";
    null;
    r2790 := (r2789);
    r2791 := "1";
    null;
    r2792 := (r2791);
    r2793 := "0";
    null;
    r2794 := (r2793);
    r2795 := "0";
    null;
    r2796 := (r2795);
    r2797 := "1";
    null;
    r2798 := (r2797);
    r2799 := "0";
    null;
    r2800 := (r2799);
    r2801 := "0";
    null;
    r2802 := (r2801);
    r2803 := "1";
    null;
    r2804 := (r2803);
    r2805 := "1";
    null;
    r2806 := (r2805);
    r2807 := "0";
    null;
    r2808 := (r2807);
    r2809 := "1";
    null;
    r2810 := (r2809);
    r2811 := "1";
    null;
    r2812 := (r2811);
    r2813 := "0";
    null;
    r2814 := (r2813);
    r2815 := "1";
    null;
    r2816 := (r2815);
    r2817 := "1";
    null;
    r2818 := (r2817);
    r2819 := "0";
    null;
    r2820 := (r2819);
    r2821 := "1";
    null;
    r2822 := (r2821);
    r2823 := "0";
    null;
    r2824 := (r2823);
    r2825 := "0";
    null;
    r2826 := (r2825);
    r2827 := "1";
    null;
    r2828 := (r2827);
    r2829 := "1";
    null;
    r2830 := (r2829);
    r2831 := "1";
    null;
    r2832 := (r2831);
    r2833 := "0";
    null;
    r2834 := (r2833);
    r2835 := "0";
    null;
    r2836 := (r2835);
    r2837 := "0";
    null;
    r2838 := (r2837);
    r2839 := "0";
    null;
    r2840 := (r2839);
    r2841 := "0";
    null;
    r2842 := (r2841);
    r2843 := "1";
    null;
    r2844 := (r2843);
    r2780 := (r2782 & r2784 & r2786 & r2788 & r2790 & r2792 & r2794 & r2796 & r2798 & r2800 & r2802 & r2804 & r2806 & r2808 & r2810 & r2812 & r2814 & r2816 & r2818 & r2820 & r2822 & r2824 & r2826 & r2828 & r2830 & r2832 & r2834 & r2836 & r2838 & r2840 & r2842 & r2844);
    return r2780;
  end rewire_MetaprogrammingRW.we49b69c1_2779;
  function rewire_MetaprogrammingRW.wc19bf174_2710 return std_logic_vector
  is
    variable r2775 : std_logic_vector(0 to 0) := (others => '0');
    variable r2774 : std_logic_vector(0 to 0) := (others => '0');
    variable r2773 : std_logic_vector(0 to 0) := (others => '0');
    variable r2772 : std_logic_vector(0 to 0) := (others => '0');
    variable r2771 : std_logic_vector(0 to 0) := (others => '0');
    variable r2770 : std_logic_vector(0 to 0) := (others => '0');
    variable r2769 : std_logic_vector(0 to 0) := (others => '0');
    variable r2768 : std_logic_vector(0 to 0) := (others => '0');
    variable r2767 : std_logic_vector(0 to 0) := (others => '0');
    variable r2766 : std_logic_vector(0 to 0) := (others => '0');
    variable r2765 : std_logic_vector(0 to 0) := (others => '0');
    variable r2764 : std_logic_vector(0 to 0) := (others => '0');
    variable r2763 : std_logic_vector(0 to 0) := (others => '0');
    variable r2762 : std_logic_vector(0 to 0) := (others => '0');
    variable r2761 : std_logic_vector(0 to 0) := (others => '0');
    variable r2760 : std_logic_vector(0 to 0) := (others => '0');
    variable r2759 : std_logic_vector(0 to 0) := (others => '0');
    variable r2758 : std_logic_vector(0 to 0) := (others => '0');
    variable r2757 : std_logic_vector(0 to 0) := (others => '0');
    variable r2756 : std_logic_vector(0 to 0) := (others => '0');
    variable r2755 : std_logic_vector(0 to 0) := (others => '0');
    variable r2754 : std_logic_vector(0 to 0) := (others => '0');
    variable r2753 : std_logic_vector(0 to 0) := (others => '0');
    variable r2752 : std_logic_vector(0 to 0) := (others => '0');
    variable r2751 : std_logic_vector(0 to 0) := (others => '0');
    variable r2750 : std_logic_vector(0 to 0) := (others => '0');
    variable r2749 : std_logic_vector(0 to 0) := (others => '0');
    variable r2748 : std_logic_vector(0 to 0) := (others => '0');
    variable r2747 : std_logic_vector(0 to 0) := (others => '0');
    variable r2746 : std_logic_vector(0 to 0) := (others => '0');
    variable r2745 : std_logic_vector(0 to 0) := (others => '0');
    variable r2744 : std_logic_vector(0 to 0) := (others => '0');
    variable r2743 : std_logic_vector(0 to 0) := (others => '0');
    variable r2742 : std_logic_vector(0 to 0) := (others => '0');
    variable r2741 : std_logic_vector(0 to 0) := (others => '0');
    variable r2740 : std_logic_vector(0 to 0) := (others => '0');
    variable r2739 : std_logic_vector(0 to 0) := (others => '0');
    variable r2738 : std_logic_vector(0 to 0) := (others => '0');
    variable r2737 : std_logic_vector(0 to 0) := (others => '0');
    variable r2736 : std_logic_vector(0 to 0) := (others => '0');
    variable r2735 : std_logic_vector(0 to 0) := (others => '0');
    variable r2734 : std_logic_vector(0 to 0) := (others => '0');
    variable r2733 : std_logic_vector(0 to 0) := (others => '0');
    variable r2732 : std_logic_vector(0 to 0) := (others => '0');
    variable r2731 : std_logic_vector(0 to 0) := (others => '0');
    variable r2730 : std_logic_vector(0 to 0) := (others => '0');
    variable r2729 : std_logic_vector(0 to 0) := (others => '0');
    variable r2728 : std_logic_vector(0 to 0) := (others => '0');
    variable r2727 : std_logic_vector(0 to 0) := (others => '0');
    variable r2726 : std_logic_vector(0 to 0) := (others => '0');
    variable r2725 : std_logic_vector(0 to 0) := (others => '0');
    variable r2724 : std_logic_vector(0 to 0) := (others => '0');
    variable r2723 : std_logic_vector(0 to 0) := (others => '0');
    variable r2722 : std_logic_vector(0 to 0) := (others => '0');
    variable r2721 : std_logic_vector(0 to 0) := (others => '0');
    variable r2720 : std_logic_vector(0 to 0) := (others => '0');
    variable r2719 : std_logic_vector(0 to 0) := (others => '0');
    variable r2718 : std_logic_vector(0 to 0) := (others => '0');
    variable r2717 : std_logic_vector(0 to 0) := (others => '0');
    variable r2716 : std_logic_vector(0 to 0) := (others => '0');
    variable r2715 : std_logic_vector(0 to 0) := (others => '0');
    variable r2714 : std_logic_vector(0 to 0) := (others => '0');
    variable r2713 : std_logic_vector(0 to 0) := (others => '0');
    variable r2712 : std_logic_vector(0 to 0) := (others => '0');
    variable r2711 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r2712 := "1";
    null;
    r2713 := (r2712);
    r2714 := "1";
    null;
    r2715 := (r2714);
    r2716 := "0";
    null;
    r2717 := (r2716);
    r2718 := "0";
    null;
    r2719 := (r2718);
    r2720 := "0";
    null;
    r2721 := (r2720);
    r2722 := "0";
    null;
    r2723 := (r2722);
    r2724 := "0";
    null;
    r2725 := (r2724);
    r2726 := "1";
    null;
    r2727 := (r2726);
    r2728 := "1";
    null;
    r2729 := (r2728);
    r2730 := "0";
    null;
    r2731 := (r2730);
    r2732 := "0";
    null;
    r2733 := (r2732);
    r2734 := "1";
    null;
    r2735 := (r2734);
    r2736 := "1";
    null;
    r2737 := (r2736);
    r2738 := "0";
    null;
    r2739 := (r2738);
    r2740 := "1";
    null;
    r2741 := (r2740);
    r2742 := "1";
    null;
    r2743 := (r2742);
    r2744 := "1";
    null;
    r2745 := (r2744);
    r2746 := "1";
    null;
    r2747 := (r2746);
    r2748 := "1";
    null;
    r2749 := (r2748);
    r2750 := "1";
    null;
    r2751 := (r2750);
    r2752 := "0";
    null;
    r2753 := (r2752);
    r2754 := "0";
    null;
    r2755 := (r2754);
    r2756 := "0";
    null;
    r2757 := (r2756);
    r2758 := "1";
    null;
    r2759 := (r2758);
    r2760 := "0";
    null;
    r2761 := (r2760);
    r2762 := "1";
    null;
    r2763 := (r2762);
    r2764 := "1";
    null;
    r2765 := (r2764);
    r2766 := "1";
    null;
    r2767 := (r2766);
    r2768 := "0";
    null;
    r2769 := (r2768);
    r2770 := "1";
    null;
    r2771 := (r2770);
    r2772 := "0";
    null;
    r2773 := (r2772);
    r2774 := "0";
    null;
    r2775 := (r2774);
    r2711 := (r2713 & r2715 & r2717 & r2719 & r2721 & r2723 & r2725 & r2727 & r2729 & r2731 & r2733 & r2735 & r2737 & r2739 & r2741 & r2743 & r2745 & r2747 & r2749 & r2751 & r2753 & r2755 & r2757 & r2759 & r2761 & r2763 & r2765 & r2767 & r2769 & r2771 & r2773 & r2775);
    return r2711;
  end rewire_MetaprogrammingRW.wc19bf174_2710;
  function rewire_MetaprogrammingRW.w9bdc06a7_2641 return std_logic_vector
  is
    variable r2706 : std_logic_vector(0 to 0) := (others => '0');
    variable r2705 : std_logic_vector(0 to 0) := (others => '0');
    variable r2704 : std_logic_vector(0 to 0) := (others => '0');
    variable r2703 : std_logic_vector(0 to 0) := (others => '0');
    variable r2702 : std_logic_vector(0 to 0) := (others => '0');
    variable r2701 : std_logic_vector(0 to 0) := (others => '0');
    variable r2700 : std_logic_vector(0 to 0) := (others => '0');
    variable r2699 : std_logic_vector(0 to 0) := (others => '0');
    variable r2698 : std_logic_vector(0 to 0) := (others => '0');
    variable r2697 : std_logic_vector(0 to 0) := (others => '0');
    variable r2696 : std_logic_vector(0 to 0) := (others => '0');
    variable r2695 : std_logic_vector(0 to 0) := (others => '0');
    variable r2694 : std_logic_vector(0 to 0) := (others => '0');
    variable r2693 : std_logic_vector(0 to 0) := (others => '0');
    variable r2692 : std_logic_vector(0 to 0) := (others => '0');
    variable r2691 : std_logic_vector(0 to 0) := (others => '0');
    variable r2690 : std_logic_vector(0 to 0) := (others => '0');
    variable r2689 : std_logic_vector(0 to 0) := (others => '0');
    variable r2688 : std_logic_vector(0 to 0) := (others => '0');
    variable r2687 : std_logic_vector(0 to 0) := (others => '0');
    variable r2686 : std_logic_vector(0 to 0) := (others => '0');
    variable r2685 : std_logic_vector(0 to 0) := (others => '0');
    variable r2684 : std_logic_vector(0 to 0) := (others => '0');
    variable r2683 : std_logic_vector(0 to 0) := (others => '0');
    variable r2682 : std_logic_vector(0 to 0) := (others => '0');
    variable r2681 : std_logic_vector(0 to 0) := (others => '0');
    variable r2680 : std_logic_vector(0 to 0) := (others => '0');
    variable r2679 : std_logic_vector(0 to 0) := (others => '0');
    variable r2678 : std_logic_vector(0 to 0) := (others => '0');
    variable r2677 : std_logic_vector(0 to 0) := (others => '0');
    variable r2676 : std_logic_vector(0 to 0) := (others => '0');
    variable r2675 : std_logic_vector(0 to 0) := (others => '0');
    variable r2674 : std_logic_vector(0 to 0) := (others => '0');
    variable r2673 : std_logic_vector(0 to 0) := (others => '0');
    variable r2672 : std_logic_vector(0 to 0) := (others => '0');
    variable r2671 : std_logic_vector(0 to 0) := (others => '0');
    variable r2670 : std_logic_vector(0 to 0) := (others => '0');
    variable r2669 : std_logic_vector(0 to 0) := (others => '0');
    variable r2668 : std_logic_vector(0 to 0) := (others => '0');
    variable r2667 : std_logic_vector(0 to 0) := (others => '0');
    variable r2666 : std_logic_vector(0 to 0) := (others => '0');
    variable r2665 : std_logic_vector(0 to 0) := (others => '0');
    variable r2664 : std_logic_vector(0 to 0) := (others => '0');
    variable r2663 : std_logic_vector(0 to 0) := (others => '0');
    variable r2662 : std_logic_vector(0 to 0) := (others => '0');
    variable r2661 : std_logic_vector(0 to 0) := (others => '0');
    variable r2660 : std_logic_vector(0 to 0) := (others => '0');
    variable r2659 : std_logic_vector(0 to 0) := (others => '0');
    variable r2658 : std_logic_vector(0 to 0) := (others => '0');
    variable r2657 : std_logic_vector(0 to 0) := (others => '0');
    variable r2656 : std_logic_vector(0 to 0) := (others => '0');
    variable r2655 : std_logic_vector(0 to 0) := (others => '0');
    variable r2654 : std_logic_vector(0 to 0) := (others => '0');
    variable r2653 : std_logic_vector(0 to 0) := (others => '0');
    variable r2652 : std_logic_vector(0 to 0) := (others => '0');
    variable r2651 : std_logic_vector(0 to 0) := (others => '0');
    variable r2650 : std_logic_vector(0 to 0) := (others => '0');
    variable r2649 : std_logic_vector(0 to 0) := (others => '0');
    variable r2648 : std_logic_vector(0 to 0) := (others => '0');
    variable r2647 : std_logic_vector(0 to 0) := (others => '0');
    variable r2646 : std_logic_vector(0 to 0) := (others => '0');
    variable r2645 : std_logic_vector(0 to 0) := (others => '0');
    variable r2644 : std_logic_vector(0 to 0) := (others => '0');
    variable r2643 : std_logic_vector(0 to 0) := (others => '0');
    variable r2642 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r2643 := "1";
    null;
    r2644 := (r2643);
    r2645 := "0";
    null;
    r2646 := (r2645);
    r2647 := "0";
    null;
    r2648 := (r2647);
    r2649 := "1";
    null;
    r2650 := (r2649);
    r2651 := "1";
    null;
    r2652 := (r2651);
    r2653 := "0";
    null;
    r2654 := (r2653);
    r2655 := "1";
    null;
    r2656 := (r2655);
    r2657 := "1";
    null;
    r2658 := (r2657);
    r2659 := "1";
    null;
    r2660 := (r2659);
    r2661 := "1";
    null;
    r2662 := (r2661);
    r2663 := "0";
    null;
    r2664 := (r2663);
    r2665 := "1";
    null;
    r2666 := (r2665);
    r2667 := "1";
    null;
    r2668 := (r2667);
    r2669 := "1";
    null;
    r2670 := (r2669);
    r2671 := "0";
    null;
    r2672 := (r2671);
    r2673 := "0";
    null;
    r2674 := (r2673);
    r2675 := "0";
    null;
    r2676 := (r2675);
    r2677 := "0";
    null;
    r2678 := (r2677);
    r2679 := "0";
    null;
    r2680 := (r2679);
    r2681 := "0";
    null;
    r2682 := (r2681);
    r2683 := "0";
    null;
    r2684 := (r2683);
    r2685 := "1";
    null;
    r2686 := (r2685);
    r2687 := "1";
    null;
    r2688 := (r2687);
    r2689 := "0";
    null;
    r2690 := (r2689);
    r2691 := "1";
    null;
    r2692 := (r2691);
    r2693 := "0";
    null;
    r2694 := (r2693);
    r2695 := "1";
    null;
    r2696 := (r2695);
    r2697 := "0";
    null;
    r2698 := (r2697);
    r2699 := "0";
    null;
    r2700 := (r2699);
    r2701 := "1";
    null;
    r2702 := (r2701);
    r2703 := "1";
    null;
    r2704 := (r2703);
    r2705 := "1";
    null;
    r2706 := (r2705);
    r2642 := (r2644 & r2646 & r2648 & r2650 & r2652 & r2654 & r2656 & r2658 & r2660 & r2662 & r2664 & r2666 & r2668 & r2670 & r2672 & r2674 & r2676 & r2678 & r2680 & r2682 & r2684 & r2686 & r2688 & r2690 & r2692 & r2694 & r2696 & r2698 & r2700 & r2702 & r2704 & r2706);
    return r2642;
  end rewire_MetaprogrammingRW.w9bdc06a7_2641;
  function rewire_MetaprogrammingRW.w80deb1fe_2572 return std_logic_vector
  is
    variable r2637 : std_logic_vector(0 to 0) := (others => '0');
    variable r2636 : std_logic_vector(0 to 0) := (others => '0');
    variable r2635 : std_logic_vector(0 to 0) := (others => '0');
    variable r2634 : std_logic_vector(0 to 0) := (others => '0');
    variable r2633 : std_logic_vector(0 to 0) := (others => '0');
    variable r2632 : std_logic_vector(0 to 0) := (others => '0');
    variable r2631 : std_logic_vector(0 to 0) := (others => '0');
    variable r2630 : std_logic_vector(0 to 0) := (others => '0');
    variable r2629 : std_logic_vector(0 to 0) := (others => '0');
    variable r2628 : std_logic_vector(0 to 0) := (others => '0');
    variable r2627 : std_logic_vector(0 to 0) := (others => '0');
    variable r2626 : std_logic_vector(0 to 0) := (others => '0');
    variable r2625 : std_logic_vector(0 to 0) := (others => '0');
    variable r2624 : std_logic_vector(0 to 0) := (others => '0');
    variable r2623 : std_logic_vector(0 to 0) := (others => '0');
    variable r2622 : std_logic_vector(0 to 0) := (others => '0');
    variable r2621 : std_logic_vector(0 to 0) := (others => '0');
    variable r2620 : std_logic_vector(0 to 0) := (others => '0');
    variable r2619 : std_logic_vector(0 to 0) := (others => '0');
    variable r2618 : std_logic_vector(0 to 0) := (others => '0');
    variable r2617 : std_logic_vector(0 to 0) := (others => '0');
    variable r2616 : std_logic_vector(0 to 0) := (others => '0');
    variable r2615 : std_logic_vector(0 to 0) := (others => '0');
    variable r2614 : std_logic_vector(0 to 0) := (others => '0');
    variable r2613 : std_logic_vector(0 to 0) := (others => '0');
    variable r2612 : std_logic_vector(0 to 0) := (others => '0');
    variable r2611 : std_logic_vector(0 to 0) := (others => '0');
    variable r2610 : std_logic_vector(0 to 0) := (others => '0');
    variable r2609 : std_logic_vector(0 to 0) := (others => '0');
    variable r2608 : std_logic_vector(0 to 0) := (others => '0');
    variable r2607 : std_logic_vector(0 to 0) := (others => '0');
    variable r2606 : std_logic_vector(0 to 0) := (others => '0');
    variable r2605 : std_logic_vector(0 to 0) := (others => '0');
    variable r2604 : std_logic_vector(0 to 0) := (others => '0');
    variable r2603 : std_logic_vector(0 to 0) := (others => '0');
    variable r2602 : std_logic_vector(0 to 0) := (others => '0');
    variable r2601 : std_logic_vector(0 to 0) := (others => '0');
    variable r2600 : std_logic_vector(0 to 0) := (others => '0');
    variable r2599 : std_logic_vector(0 to 0) := (others => '0');
    variable r2598 : std_logic_vector(0 to 0) := (others => '0');
    variable r2597 : std_logic_vector(0 to 0) := (others => '0');
    variable r2596 : std_logic_vector(0 to 0) := (others => '0');
    variable r2595 : std_logic_vector(0 to 0) := (others => '0');
    variable r2594 : std_logic_vector(0 to 0) := (others => '0');
    variable r2593 : std_logic_vector(0 to 0) := (others => '0');
    variable r2592 : std_logic_vector(0 to 0) := (others => '0');
    variable r2591 : std_logic_vector(0 to 0) := (others => '0');
    variable r2590 : std_logic_vector(0 to 0) := (others => '0');
    variable r2589 : std_logic_vector(0 to 0) := (others => '0');
    variable r2588 : std_logic_vector(0 to 0) := (others => '0');
    variable r2587 : std_logic_vector(0 to 0) := (others => '0');
    variable r2586 : std_logic_vector(0 to 0) := (others => '0');
    variable r2585 : std_logic_vector(0 to 0) := (others => '0');
    variable r2584 : std_logic_vector(0 to 0) := (others => '0');
    variable r2583 : std_logic_vector(0 to 0) := (others => '0');
    variable r2582 : std_logic_vector(0 to 0) := (others => '0');
    variable r2581 : std_logic_vector(0 to 0) := (others => '0');
    variable r2580 : std_logic_vector(0 to 0) := (others => '0');
    variable r2579 : std_logic_vector(0 to 0) := (others => '0');
    variable r2578 : std_logic_vector(0 to 0) := (others => '0');
    variable r2577 : std_logic_vector(0 to 0) := (others => '0');
    variable r2576 : std_logic_vector(0 to 0) := (others => '0');
    variable r2575 : std_logic_vector(0 to 0) := (others => '0');
    variable r2574 : std_logic_vector(0 to 0) := (others => '0');
    variable r2573 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r2574 := "1";
    null;
    r2575 := (r2574);
    r2576 := "0";
    null;
    r2577 := (r2576);
    r2578 := "0";
    null;
    r2579 := (r2578);
    r2580 := "0";
    null;
    r2581 := (r2580);
    r2582 := "0";
    null;
    r2583 := (r2582);
    r2584 := "0";
    null;
    r2585 := (r2584);
    r2586 := "0";
    null;
    r2587 := (r2586);
    r2588 := "0";
    null;
    r2589 := (r2588);
    r2590 := "1";
    null;
    r2591 := (r2590);
    r2592 := "1";
    null;
    r2593 := (r2592);
    r2594 := "0";
    null;
    r2595 := (r2594);
    r2596 := "1";
    null;
    r2597 := (r2596);
    r2598 := "1";
    null;
    r2599 := (r2598);
    r2600 := "1";
    null;
    r2601 := (r2600);
    r2602 := "1";
    null;
    r2603 := (r2602);
    r2604 := "0";
    null;
    r2605 := (r2604);
    r2606 := "1";
    null;
    r2607 := (r2606);
    r2608 := "0";
    null;
    r2609 := (r2608);
    r2610 := "1";
    null;
    r2611 := (r2610);
    r2612 := "1";
    null;
    r2613 := (r2612);
    r2614 := "0";
    null;
    r2615 := (r2614);
    r2616 := "0";
    null;
    r2617 := (r2616);
    r2618 := "0";
    null;
    r2619 := (r2618);
    r2620 := "1";
    null;
    r2621 := (r2620);
    r2622 := "1";
    null;
    r2623 := (r2622);
    r2624 := "1";
    null;
    r2625 := (r2624);
    r2626 := "1";
    null;
    r2627 := (r2626);
    r2628 := "1";
    null;
    r2629 := (r2628);
    r2630 := "1";
    null;
    r2631 := (r2630);
    r2632 := "1";
    null;
    r2633 := (r2632);
    r2634 := "1";
    null;
    r2635 := (r2634);
    r2636 := "0";
    null;
    r2637 := (r2636);
    r2573 := (r2575 & r2577 & r2579 & r2581 & r2583 & r2585 & r2587 & r2589 & r2591 & r2593 & r2595 & r2597 & r2599 & r2601 & r2603 & r2605 & r2607 & r2609 & r2611 & r2613 & r2615 & r2617 & r2619 & r2621 & r2623 & r2625 & r2627 & r2629 & r2631 & r2633 & r2635 & r2637);
    return r2573;
  end rewire_MetaprogrammingRW.w80deb1fe_2572;
  function rewire_MetaprogrammingRW.w72be5d74_2503 return std_logic_vector
  is
    variable r2568 : std_logic_vector(0 to 0) := (others => '0');
    variable r2567 : std_logic_vector(0 to 0) := (others => '0');
    variable r2566 : std_logic_vector(0 to 0) := (others => '0');
    variable r2565 : std_logic_vector(0 to 0) := (others => '0');
    variable r2564 : std_logic_vector(0 to 0) := (others => '0');
    variable r2563 : std_logic_vector(0 to 0) := (others => '0');
    variable r2562 : std_logic_vector(0 to 0) := (others => '0');
    variable r2561 : std_logic_vector(0 to 0) := (others => '0');
    variable r2560 : std_logic_vector(0 to 0) := (others => '0');
    variable r2559 : std_logic_vector(0 to 0) := (others => '0');
    variable r2558 : std_logic_vector(0 to 0) := (others => '0');
    variable r2557 : std_logic_vector(0 to 0) := (others => '0');
    variable r2556 : std_logic_vector(0 to 0) := (others => '0');
    variable r2555 : std_logic_vector(0 to 0) := (others => '0');
    variable r2554 : std_logic_vector(0 to 0) := (others => '0');
    variable r2553 : std_logic_vector(0 to 0) := (others => '0');
    variable r2552 : std_logic_vector(0 to 0) := (others => '0');
    variable r2551 : std_logic_vector(0 to 0) := (others => '0');
    variable r2550 : std_logic_vector(0 to 0) := (others => '0');
    variable r2549 : std_logic_vector(0 to 0) := (others => '0');
    variable r2548 : std_logic_vector(0 to 0) := (others => '0');
    variable r2547 : std_logic_vector(0 to 0) := (others => '0');
    variable r2546 : std_logic_vector(0 to 0) := (others => '0');
    variable r2545 : std_logic_vector(0 to 0) := (others => '0');
    variable r2544 : std_logic_vector(0 to 0) := (others => '0');
    variable r2543 : std_logic_vector(0 to 0) := (others => '0');
    variable r2542 : std_logic_vector(0 to 0) := (others => '0');
    variable r2541 : std_logic_vector(0 to 0) := (others => '0');
    variable r2540 : std_logic_vector(0 to 0) := (others => '0');
    variable r2539 : std_logic_vector(0 to 0) := (others => '0');
    variable r2538 : std_logic_vector(0 to 0) := (others => '0');
    variable r2537 : std_logic_vector(0 to 0) := (others => '0');
    variable r2536 : std_logic_vector(0 to 0) := (others => '0');
    variable r2535 : std_logic_vector(0 to 0) := (others => '0');
    variable r2534 : std_logic_vector(0 to 0) := (others => '0');
    variable r2533 : std_logic_vector(0 to 0) := (others => '0');
    variable r2532 : std_logic_vector(0 to 0) := (others => '0');
    variable r2531 : std_logic_vector(0 to 0) := (others => '0');
    variable r2530 : std_logic_vector(0 to 0) := (others => '0');
    variable r2529 : std_logic_vector(0 to 0) := (others => '0');
    variable r2528 : std_logic_vector(0 to 0) := (others => '0');
    variable r2527 : std_logic_vector(0 to 0) := (others => '0');
    variable r2526 : std_logic_vector(0 to 0) := (others => '0');
    variable r2525 : std_logic_vector(0 to 0) := (others => '0');
    variable r2524 : std_logic_vector(0 to 0) := (others => '0');
    variable r2523 : std_logic_vector(0 to 0) := (others => '0');
    variable r2522 : std_logic_vector(0 to 0) := (others => '0');
    variable r2521 : std_logic_vector(0 to 0) := (others => '0');
    variable r2520 : std_logic_vector(0 to 0) := (others => '0');
    variable r2519 : std_logic_vector(0 to 0) := (others => '0');
    variable r2518 : std_logic_vector(0 to 0) := (others => '0');
    variable r2517 : std_logic_vector(0 to 0) := (others => '0');
    variable r2516 : std_logic_vector(0 to 0) := (others => '0');
    variable r2515 : std_logic_vector(0 to 0) := (others => '0');
    variable r2514 : std_logic_vector(0 to 0) := (others => '0');
    variable r2513 : std_logic_vector(0 to 0) := (others => '0');
    variable r2512 : std_logic_vector(0 to 0) := (others => '0');
    variable r2511 : std_logic_vector(0 to 0) := (others => '0');
    variable r2510 : std_logic_vector(0 to 0) := (others => '0');
    variable r2509 : std_logic_vector(0 to 0) := (others => '0');
    variable r2508 : std_logic_vector(0 to 0) := (others => '0');
    variable r2507 : std_logic_vector(0 to 0) := (others => '0');
    variable r2506 : std_logic_vector(0 to 0) := (others => '0');
    variable r2505 : std_logic_vector(0 to 0) := (others => '0');
    variable r2504 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r2505 := "0";
    null;
    r2506 := (r2505);
    r2507 := "1";
    null;
    r2508 := (r2507);
    r2509 := "1";
    null;
    r2510 := (r2509);
    r2511 := "1";
    null;
    r2512 := (r2511);
    r2513 := "0";
    null;
    r2514 := (r2513);
    r2515 := "0";
    null;
    r2516 := (r2515);
    r2517 := "1";
    null;
    r2518 := (r2517);
    r2519 := "0";
    null;
    r2520 := (r2519);
    r2521 := "1";
    null;
    r2522 := (r2521);
    r2523 := "0";
    null;
    r2524 := (r2523);
    r2525 := "1";
    null;
    r2526 := (r2525);
    r2527 := "1";
    null;
    r2528 := (r2527);
    r2529 := "1";
    null;
    r2530 := (r2529);
    r2531 := "1";
    null;
    r2532 := (r2531);
    r2533 := "1";
    null;
    r2534 := (r2533);
    r2535 := "0";
    null;
    r2536 := (r2535);
    r2537 := "0";
    null;
    r2538 := (r2537);
    r2539 := "1";
    null;
    r2540 := (r2539);
    r2541 := "0";
    null;
    r2542 := (r2541);
    r2543 := "1";
    null;
    r2544 := (r2543);
    r2545 := "1";
    null;
    r2546 := (r2545);
    r2547 := "1";
    null;
    r2548 := (r2547);
    r2549 := "0";
    null;
    r2550 := (r2549);
    r2551 := "1";
    null;
    r2552 := (r2551);
    r2553 := "0";
    null;
    r2554 := (r2553);
    r2555 := "1";
    null;
    r2556 := (r2555);
    r2557 := "1";
    null;
    r2558 := (r2557);
    r2559 := "1";
    null;
    r2560 := (r2559);
    r2561 := "0";
    null;
    r2562 := (r2561);
    r2563 := "1";
    null;
    r2564 := (r2563);
    r2565 := "0";
    null;
    r2566 := (r2565);
    r2567 := "0";
    null;
    r2568 := (r2567);
    r2504 := (r2506 & r2508 & r2510 & r2512 & r2514 & r2516 & r2518 & r2520 & r2522 & r2524 & r2526 & r2528 & r2530 & r2532 & r2534 & r2536 & r2538 & r2540 & r2542 & r2544 & r2546 & r2548 & r2550 & r2552 & r2554 & r2556 & r2558 & r2560 & r2562 & r2564 & r2566 & r2568);
    return r2504;
  end rewire_MetaprogrammingRW.w72be5d74_2503;
  function rewire_MetaprogrammingRW.w550c7dc3_2434 return std_logic_vector
  is
    variable r2499 : std_logic_vector(0 to 0) := (others => '0');
    variable r2498 : std_logic_vector(0 to 0) := (others => '0');
    variable r2497 : std_logic_vector(0 to 0) := (others => '0');
    variable r2496 : std_logic_vector(0 to 0) := (others => '0');
    variable r2495 : std_logic_vector(0 to 0) := (others => '0');
    variable r2494 : std_logic_vector(0 to 0) := (others => '0');
    variable r2493 : std_logic_vector(0 to 0) := (others => '0');
    variable r2492 : std_logic_vector(0 to 0) := (others => '0');
    variable r2491 : std_logic_vector(0 to 0) := (others => '0');
    variable r2490 : std_logic_vector(0 to 0) := (others => '0');
    variable r2489 : std_logic_vector(0 to 0) := (others => '0');
    variable r2488 : std_logic_vector(0 to 0) := (others => '0');
    variable r2487 : std_logic_vector(0 to 0) := (others => '0');
    variable r2486 : std_logic_vector(0 to 0) := (others => '0');
    variable r2485 : std_logic_vector(0 to 0) := (others => '0');
    variable r2484 : std_logic_vector(0 to 0) := (others => '0');
    variable r2483 : std_logic_vector(0 to 0) := (others => '0');
    variable r2482 : std_logic_vector(0 to 0) := (others => '0');
    variable r2481 : std_logic_vector(0 to 0) := (others => '0');
    variable r2480 : std_logic_vector(0 to 0) := (others => '0');
    variable r2479 : std_logic_vector(0 to 0) := (others => '0');
    variable r2478 : std_logic_vector(0 to 0) := (others => '0');
    variable r2477 : std_logic_vector(0 to 0) := (others => '0');
    variable r2476 : std_logic_vector(0 to 0) := (others => '0');
    variable r2475 : std_logic_vector(0 to 0) := (others => '0');
    variable r2474 : std_logic_vector(0 to 0) := (others => '0');
    variable r2473 : std_logic_vector(0 to 0) := (others => '0');
    variable r2472 : std_logic_vector(0 to 0) := (others => '0');
    variable r2471 : std_logic_vector(0 to 0) := (others => '0');
    variable r2470 : std_logic_vector(0 to 0) := (others => '0');
    variable r2469 : std_logic_vector(0 to 0) := (others => '0');
    variable r2468 : std_logic_vector(0 to 0) := (others => '0');
    variable r2467 : std_logic_vector(0 to 0) := (others => '0');
    variable r2466 : std_logic_vector(0 to 0) := (others => '0');
    variable r2465 : std_logic_vector(0 to 0) := (others => '0');
    variable r2464 : std_logic_vector(0 to 0) := (others => '0');
    variable r2463 : std_logic_vector(0 to 0) := (others => '0');
    variable r2462 : std_logic_vector(0 to 0) := (others => '0');
    variable r2461 : std_logic_vector(0 to 0) := (others => '0');
    variable r2460 : std_logic_vector(0 to 0) := (others => '0');
    variable r2459 : std_logic_vector(0 to 0) := (others => '0');
    variable r2458 : std_logic_vector(0 to 0) := (others => '0');
    variable r2457 : std_logic_vector(0 to 0) := (others => '0');
    variable r2456 : std_logic_vector(0 to 0) := (others => '0');
    variable r2455 : std_logic_vector(0 to 0) := (others => '0');
    variable r2454 : std_logic_vector(0 to 0) := (others => '0');
    variable r2453 : std_logic_vector(0 to 0) := (others => '0');
    variable r2452 : std_logic_vector(0 to 0) := (others => '0');
    variable r2451 : std_logic_vector(0 to 0) := (others => '0');
    variable r2450 : std_logic_vector(0 to 0) := (others => '0');
    variable r2449 : std_logic_vector(0 to 0) := (others => '0');
    variable r2448 : std_logic_vector(0 to 0) := (others => '0');
    variable r2447 : std_logic_vector(0 to 0) := (others => '0');
    variable r2446 : std_logic_vector(0 to 0) := (others => '0');
    variable r2445 : std_logic_vector(0 to 0) := (others => '0');
    variable r2444 : std_logic_vector(0 to 0) := (others => '0');
    variable r2443 : std_logic_vector(0 to 0) := (others => '0');
    variable r2442 : std_logic_vector(0 to 0) := (others => '0');
    variable r2441 : std_logic_vector(0 to 0) := (others => '0');
    variable r2440 : std_logic_vector(0 to 0) := (others => '0');
    variable r2439 : std_logic_vector(0 to 0) := (others => '0');
    variable r2438 : std_logic_vector(0 to 0) := (others => '0');
    variable r2437 : std_logic_vector(0 to 0) := (others => '0');
    variable r2436 : std_logic_vector(0 to 0) := (others => '0');
    variable r2435 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r2436 := "0";
    null;
    r2437 := (r2436);
    r2438 := "1";
    null;
    r2439 := (r2438);
    r2440 := "0";
    null;
    r2441 := (r2440);
    r2442 := "1";
    null;
    r2443 := (r2442);
    r2444 := "0";
    null;
    r2445 := (r2444);
    r2446 := "1";
    null;
    r2447 := (r2446);
    r2448 := "0";
    null;
    r2449 := (r2448);
    r2450 := "1";
    null;
    r2451 := (r2450);
    r2452 := "0";
    null;
    r2453 := (r2452);
    r2454 := "0";
    null;
    r2455 := (r2454);
    r2456 := "0";
    null;
    r2457 := (r2456);
    r2458 := "0";
    null;
    r2459 := (r2458);
    r2460 := "1";
    null;
    r2461 := (r2460);
    r2462 := "1";
    null;
    r2463 := (r2462);
    r2464 := "0";
    null;
    r2465 := (r2464);
    r2466 := "0";
    null;
    r2467 := (r2466);
    r2468 := "0";
    null;
    r2469 := (r2468);
    r2470 := "1";
    null;
    r2471 := (r2470);
    r2472 := "1";
    null;
    r2473 := (r2472);
    r2474 := "1";
    null;
    r2475 := (r2474);
    r2476 := "1";
    null;
    r2477 := (r2476);
    r2478 := "1";
    null;
    r2479 := (r2478);
    r2480 := "0";
    null;
    r2481 := (r2480);
    r2482 := "1";
    null;
    r2483 := (r2482);
    r2484 := "1";
    null;
    r2485 := (r2484);
    r2486 := "1";
    null;
    r2487 := (r2486);
    r2488 := "0";
    null;
    r2489 := (r2488);
    r2490 := "0";
    null;
    r2491 := (r2490);
    r2492 := "0";
    null;
    r2493 := (r2492);
    r2494 := "0";
    null;
    r2495 := (r2494);
    r2496 := "1";
    null;
    r2497 := (r2496);
    r2498 := "1";
    null;
    r2499 := (r2498);
    r2435 := (r2437 & r2439 & r2441 & r2443 & r2445 & r2447 & r2449 & r2451 & r2453 & r2455 & r2457 & r2459 & r2461 & r2463 & r2465 & r2467 & r2469 & r2471 & r2473 & r2475 & r2477 & r2479 & r2481 & r2483 & r2485 & r2487 & r2489 & r2491 & r2493 & r2495 & r2497 & r2499);
    return r2435;
  end rewire_MetaprogrammingRW.w550c7dc3_2434;
  function rewire_MetaprogrammingRW.w243185be_2365 return std_logic_vector
  is
    variable r2430 : std_logic_vector(0 to 0) := (others => '0');
    variable r2429 : std_logic_vector(0 to 0) := (others => '0');
    variable r2428 : std_logic_vector(0 to 0) := (others => '0');
    variable r2427 : std_logic_vector(0 to 0) := (others => '0');
    variable r2426 : std_logic_vector(0 to 0) := (others => '0');
    variable r2425 : std_logic_vector(0 to 0) := (others => '0');
    variable r2424 : std_logic_vector(0 to 0) := (others => '0');
    variable r2423 : std_logic_vector(0 to 0) := (others => '0');
    variable r2422 : std_logic_vector(0 to 0) := (others => '0');
    variable r2421 : std_logic_vector(0 to 0) := (others => '0');
    variable r2420 : std_logic_vector(0 to 0) := (others => '0');
    variable r2419 : std_logic_vector(0 to 0) := (others => '0');
    variable r2418 : std_logic_vector(0 to 0) := (others => '0');
    variable r2417 : std_logic_vector(0 to 0) := (others => '0');
    variable r2416 : std_logic_vector(0 to 0) := (others => '0');
    variable r2415 : std_logic_vector(0 to 0) := (others => '0');
    variable r2414 : std_logic_vector(0 to 0) := (others => '0');
    variable r2413 : std_logic_vector(0 to 0) := (others => '0');
    variable r2412 : std_logic_vector(0 to 0) := (others => '0');
    variable r2411 : std_logic_vector(0 to 0) := (others => '0');
    variable r2410 : std_logic_vector(0 to 0) := (others => '0');
    variable r2409 : std_logic_vector(0 to 0) := (others => '0');
    variable r2408 : std_logic_vector(0 to 0) := (others => '0');
    variable r2407 : std_logic_vector(0 to 0) := (others => '0');
    variable r2406 : std_logic_vector(0 to 0) := (others => '0');
    variable r2405 : std_logic_vector(0 to 0) := (others => '0');
    variable r2404 : std_logic_vector(0 to 0) := (others => '0');
    variable r2403 : std_logic_vector(0 to 0) := (others => '0');
    variable r2402 : std_logic_vector(0 to 0) := (others => '0');
    variable r2401 : std_logic_vector(0 to 0) := (others => '0');
    variable r2400 : std_logic_vector(0 to 0) := (others => '0');
    variable r2399 : std_logic_vector(0 to 0) := (others => '0');
    variable r2398 : std_logic_vector(0 to 0) := (others => '0');
    variable r2397 : std_logic_vector(0 to 0) := (others => '0');
    variable r2396 : std_logic_vector(0 to 0) := (others => '0');
    variable r2395 : std_logic_vector(0 to 0) := (others => '0');
    variable r2394 : std_logic_vector(0 to 0) := (others => '0');
    variable r2393 : std_logic_vector(0 to 0) := (others => '0');
    variable r2392 : std_logic_vector(0 to 0) := (others => '0');
    variable r2391 : std_logic_vector(0 to 0) := (others => '0');
    variable r2390 : std_logic_vector(0 to 0) := (others => '0');
    variable r2389 : std_logic_vector(0 to 0) := (others => '0');
    variable r2388 : std_logic_vector(0 to 0) := (others => '0');
    variable r2387 : std_logic_vector(0 to 0) := (others => '0');
    variable r2386 : std_logic_vector(0 to 0) := (others => '0');
    variable r2385 : std_logic_vector(0 to 0) := (others => '0');
    variable r2384 : std_logic_vector(0 to 0) := (others => '0');
    variable r2383 : std_logic_vector(0 to 0) := (others => '0');
    variable r2382 : std_logic_vector(0 to 0) := (others => '0');
    variable r2381 : std_logic_vector(0 to 0) := (others => '0');
    variable r2380 : std_logic_vector(0 to 0) := (others => '0');
    variable r2379 : std_logic_vector(0 to 0) := (others => '0');
    variable r2378 : std_logic_vector(0 to 0) := (others => '0');
    variable r2377 : std_logic_vector(0 to 0) := (others => '0');
    variable r2376 : std_logic_vector(0 to 0) := (others => '0');
    variable r2375 : std_logic_vector(0 to 0) := (others => '0');
    variable r2374 : std_logic_vector(0 to 0) := (others => '0');
    variable r2373 : std_logic_vector(0 to 0) := (others => '0');
    variable r2372 : std_logic_vector(0 to 0) := (others => '0');
    variable r2371 : std_logic_vector(0 to 0) := (others => '0');
    variable r2370 : std_logic_vector(0 to 0) := (others => '0');
    variable r2369 : std_logic_vector(0 to 0) := (others => '0');
    variable r2368 : std_logic_vector(0 to 0) := (others => '0');
    variable r2367 : std_logic_vector(0 to 0) := (others => '0');
    variable r2366 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r2367 := "0";
    null;
    r2368 := (r2367);
    r2369 := "0";
    null;
    r2370 := (r2369);
    r2371 := "1";
    null;
    r2372 := (r2371);
    r2373 := "0";
    null;
    r2374 := (r2373);
    r2375 := "0";
    null;
    r2376 := (r2375);
    r2377 := "1";
    null;
    r2378 := (r2377);
    r2379 := "0";
    null;
    r2380 := (r2379);
    r2381 := "0";
    null;
    r2382 := (r2381);
    r2383 := "0";
    null;
    r2384 := (r2383);
    r2385 := "0";
    null;
    r2386 := (r2385);
    r2387 := "1";
    null;
    r2388 := (r2387);
    r2389 := "1";
    null;
    r2390 := (r2389);
    r2391 := "0";
    null;
    r2392 := (r2391);
    r2393 := "0";
    null;
    r2394 := (r2393);
    r2395 := "0";
    null;
    r2396 := (r2395);
    r2397 := "1";
    null;
    r2398 := (r2397);
    r2399 := "1";
    null;
    r2400 := (r2399);
    r2401 := "0";
    null;
    r2402 := (r2401);
    r2403 := "0";
    null;
    r2404 := (r2403);
    r2405 := "0";
    null;
    r2406 := (r2405);
    r2407 := "0";
    null;
    r2408 := (r2407);
    r2409 := "1";
    null;
    r2410 := (r2409);
    r2411 := "0";
    null;
    r2412 := (r2411);
    r2413 := "1";
    null;
    r2414 := (r2413);
    r2415 := "1";
    null;
    r2416 := (r2415);
    r2417 := "0";
    null;
    r2418 := (r2417);
    r2419 := "1";
    null;
    r2420 := (r2419);
    r2421 := "1";
    null;
    r2422 := (r2421);
    r2423 := "1";
    null;
    r2424 := (r2423);
    r2425 := "1";
    null;
    r2426 := (r2425);
    r2427 := "1";
    null;
    r2428 := (r2427);
    r2429 := "0";
    null;
    r2430 := (r2429);
    r2366 := (r2368 & r2370 & r2372 & r2374 & r2376 & r2378 & r2380 & r2382 & r2384 & r2386 & r2388 & r2390 & r2392 & r2394 & r2396 & r2398 & r2400 & r2402 & r2404 & r2406 & r2408 & r2410 & r2412 & r2414 & r2416 & r2418 & r2420 & r2422 & r2424 & r2426 & r2428 & r2430);
    return r2366;
  end rewire_MetaprogrammingRW.w243185be_2365;
  function rewire_MetaprogrammingRW.w12835b01_2296 return std_logic_vector
  is
    variable r2361 : std_logic_vector(0 to 0) := (others => '0');
    variable r2360 : std_logic_vector(0 to 0) := (others => '0');
    variable r2359 : std_logic_vector(0 to 0) := (others => '0');
    variable r2358 : std_logic_vector(0 to 0) := (others => '0');
    variable r2357 : std_logic_vector(0 to 0) := (others => '0');
    variable r2356 : std_logic_vector(0 to 0) := (others => '0');
    variable r2355 : std_logic_vector(0 to 0) := (others => '0');
    variable r2354 : std_logic_vector(0 to 0) := (others => '0');
    variable r2353 : std_logic_vector(0 to 0) := (others => '0');
    variable r2352 : std_logic_vector(0 to 0) := (others => '0');
    variable r2351 : std_logic_vector(0 to 0) := (others => '0');
    variable r2350 : std_logic_vector(0 to 0) := (others => '0');
    variable r2349 : std_logic_vector(0 to 0) := (others => '0');
    variable r2348 : std_logic_vector(0 to 0) := (others => '0');
    variable r2347 : std_logic_vector(0 to 0) := (others => '0');
    variable r2346 : std_logic_vector(0 to 0) := (others => '0');
    variable r2345 : std_logic_vector(0 to 0) := (others => '0');
    variable r2344 : std_logic_vector(0 to 0) := (others => '0');
    variable r2343 : std_logic_vector(0 to 0) := (others => '0');
    variable r2342 : std_logic_vector(0 to 0) := (others => '0');
    variable r2341 : std_logic_vector(0 to 0) := (others => '0');
    variable r2340 : std_logic_vector(0 to 0) := (others => '0');
    variable r2339 : std_logic_vector(0 to 0) := (others => '0');
    variable r2338 : std_logic_vector(0 to 0) := (others => '0');
    variable r2337 : std_logic_vector(0 to 0) := (others => '0');
    variable r2336 : std_logic_vector(0 to 0) := (others => '0');
    variable r2335 : std_logic_vector(0 to 0) := (others => '0');
    variable r2334 : std_logic_vector(0 to 0) := (others => '0');
    variable r2333 : std_logic_vector(0 to 0) := (others => '0');
    variable r2332 : std_logic_vector(0 to 0) := (others => '0');
    variable r2331 : std_logic_vector(0 to 0) := (others => '0');
    variable r2330 : std_logic_vector(0 to 0) := (others => '0');
    variable r2329 : std_logic_vector(0 to 0) := (others => '0');
    variable r2328 : std_logic_vector(0 to 0) := (others => '0');
    variable r2327 : std_logic_vector(0 to 0) := (others => '0');
    variable r2326 : std_logic_vector(0 to 0) := (others => '0');
    variable r2325 : std_logic_vector(0 to 0) := (others => '0');
    variable r2324 : std_logic_vector(0 to 0) := (others => '0');
    variable r2323 : std_logic_vector(0 to 0) := (others => '0');
    variable r2322 : std_logic_vector(0 to 0) := (others => '0');
    variable r2321 : std_logic_vector(0 to 0) := (others => '0');
    variable r2320 : std_logic_vector(0 to 0) := (others => '0');
    variable r2319 : std_logic_vector(0 to 0) := (others => '0');
    variable r2318 : std_logic_vector(0 to 0) := (others => '0');
    variable r2317 : std_logic_vector(0 to 0) := (others => '0');
    variable r2316 : std_logic_vector(0 to 0) := (others => '0');
    variable r2315 : std_logic_vector(0 to 0) := (others => '0');
    variable r2314 : std_logic_vector(0 to 0) := (others => '0');
    variable r2313 : std_logic_vector(0 to 0) := (others => '0');
    variable r2312 : std_logic_vector(0 to 0) := (others => '0');
    variable r2311 : std_logic_vector(0 to 0) := (others => '0');
    variable r2310 : std_logic_vector(0 to 0) := (others => '0');
    variable r2309 : std_logic_vector(0 to 0) := (others => '0');
    variable r2308 : std_logic_vector(0 to 0) := (others => '0');
    variable r2307 : std_logic_vector(0 to 0) := (others => '0');
    variable r2306 : std_logic_vector(0 to 0) := (others => '0');
    variable r2305 : std_logic_vector(0 to 0) := (others => '0');
    variable r2304 : std_logic_vector(0 to 0) := (others => '0');
    variable r2303 : std_logic_vector(0 to 0) := (others => '0');
    variable r2302 : std_logic_vector(0 to 0) := (others => '0');
    variable r2301 : std_logic_vector(0 to 0) := (others => '0');
    variable r2300 : std_logic_vector(0 to 0) := (others => '0');
    variable r2299 : std_logic_vector(0 to 0) := (others => '0');
    variable r2298 : std_logic_vector(0 to 0) := (others => '0');
    variable r2297 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r2298 := "0";
    null;
    r2299 := (r2298);
    r2300 := "0";
    null;
    r2301 := (r2300);
    r2302 := "0";
    null;
    r2303 := (r2302);
    r2304 := "1";
    null;
    r2305 := (r2304);
    r2306 := "0";
    null;
    r2307 := (r2306);
    r2308 := "0";
    null;
    r2309 := (r2308);
    r2310 := "1";
    null;
    r2311 := (r2310);
    r2312 := "0";
    null;
    r2313 := (r2312);
    r2314 := "1";
    null;
    r2315 := (r2314);
    r2316 := "0";
    null;
    r2317 := (r2316);
    r2318 := "0";
    null;
    r2319 := (r2318);
    r2320 := "0";
    null;
    r2321 := (r2320);
    r2322 := "0";
    null;
    r2323 := (r2322);
    r2324 := "0";
    null;
    r2325 := (r2324);
    r2326 := "1";
    null;
    r2327 := (r2326);
    r2328 := "1";
    null;
    r2329 := (r2328);
    r2330 := "0";
    null;
    r2331 := (r2330);
    r2332 := "1";
    null;
    r2333 := (r2332);
    r2334 := "0";
    null;
    r2335 := (r2334);
    r2336 := "1";
    null;
    r2337 := (r2336);
    r2338 := "1";
    null;
    r2339 := (r2338);
    r2340 := "0";
    null;
    r2341 := (r2340);
    r2342 := "1";
    null;
    r2343 := (r2342);
    r2344 := "1";
    null;
    r2345 := (r2344);
    r2346 := "0";
    null;
    r2347 := (r2346);
    r2348 := "0";
    null;
    r2349 := (r2348);
    r2350 := "0";
    null;
    r2351 := (r2350);
    r2352 := "0";
    null;
    r2353 := (r2352);
    r2354 := "0";
    null;
    r2355 := (r2354);
    r2356 := "0";
    null;
    r2357 := (r2356);
    r2358 := "0";
    null;
    r2359 := (r2358);
    r2360 := "1";
    null;
    r2361 := (r2360);
    r2297 := (r2299 & r2301 & r2303 & r2305 & r2307 & r2309 & r2311 & r2313 & r2315 & r2317 & r2319 & r2321 & r2323 & r2325 & r2327 & r2329 & r2331 & r2333 & r2335 & r2337 & r2339 & r2341 & r2343 & r2345 & r2347 & r2349 & r2351 & r2353 & r2355 & r2357 & r2359 & r2361);
    return r2297;
  end rewire_MetaprogrammingRW.w12835b01_2296;
  function rewire_MetaprogrammingRW.wd807aa98_2227 return std_logic_vector
  is
    variable r2292 : std_logic_vector(0 to 0) := (others => '0');
    variable r2291 : std_logic_vector(0 to 0) := (others => '0');
    variable r2290 : std_logic_vector(0 to 0) := (others => '0');
    variable r2289 : std_logic_vector(0 to 0) := (others => '0');
    variable r2288 : std_logic_vector(0 to 0) := (others => '0');
    variable r2287 : std_logic_vector(0 to 0) := (others => '0');
    variable r2286 : std_logic_vector(0 to 0) := (others => '0');
    variable r2285 : std_logic_vector(0 to 0) := (others => '0');
    variable r2284 : std_logic_vector(0 to 0) := (others => '0');
    variable r2283 : std_logic_vector(0 to 0) := (others => '0');
    variable r2282 : std_logic_vector(0 to 0) := (others => '0');
    variable r2281 : std_logic_vector(0 to 0) := (others => '0');
    variable r2280 : std_logic_vector(0 to 0) := (others => '0');
    variable r2279 : std_logic_vector(0 to 0) := (others => '0');
    variable r2278 : std_logic_vector(0 to 0) := (others => '0');
    variable r2277 : std_logic_vector(0 to 0) := (others => '0');
    variable r2276 : std_logic_vector(0 to 0) := (others => '0');
    variable r2275 : std_logic_vector(0 to 0) := (others => '0');
    variable r2274 : std_logic_vector(0 to 0) := (others => '0');
    variable r2273 : std_logic_vector(0 to 0) := (others => '0');
    variable r2272 : std_logic_vector(0 to 0) := (others => '0');
    variable r2271 : std_logic_vector(0 to 0) := (others => '0');
    variable r2270 : std_logic_vector(0 to 0) := (others => '0');
    variable r2269 : std_logic_vector(0 to 0) := (others => '0');
    variable r2268 : std_logic_vector(0 to 0) := (others => '0');
    variable r2267 : std_logic_vector(0 to 0) := (others => '0');
    variable r2266 : std_logic_vector(0 to 0) := (others => '0');
    variable r2265 : std_logic_vector(0 to 0) := (others => '0');
    variable r2264 : std_logic_vector(0 to 0) := (others => '0');
    variable r2263 : std_logic_vector(0 to 0) := (others => '0');
    variable r2262 : std_logic_vector(0 to 0) := (others => '0');
    variable r2261 : std_logic_vector(0 to 0) := (others => '0');
    variable r2260 : std_logic_vector(0 to 0) := (others => '0');
    variable r2259 : std_logic_vector(0 to 0) := (others => '0');
    variable r2258 : std_logic_vector(0 to 0) := (others => '0');
    variable r2257 : std_logic_vector(0 to 0) := (others => '0');
    variable r2256 : std_logic_vector(0 to 0) := (others => '0');
    variable r2255 : std_logic_vector(0 to 0) := (others => '0');
    variable r2254 : std_logic_vector(0 to 0) := (others => '0');
    variable r2253 : std_logic_vector(0 to 0) := (others => '0');
    variable r2252 : std_logic_vector(0 to 0) := (others => '0');
    variable r2251 : std_logic_vector(0 to 0) := (others => '0');
    variable r2250 : std_logic_vector(0 to 0) := (others => '0');
    variable r2249 : std_logic_vector(0 to 0) := (others => '0');
    variable r2248 : std_logic_vector(0 to 0) := (others => '0');
    variable r2247 : std_logic_vector(0 to 0) := (others => '0');
    variable r2246 : std_logic_vector(0 to 0) := (others => '0');
    variable r2245 : std_logic_vector(0 to 0) := (others => '0');
    variable r2244 : std_logic_vector(0 to 0) := (others => '0');
    variable r2243 : std_logic_vector(0 to 0) := (others => '0');
    variable r2242 : std_logic_vector(0 to 0) := (others => '0');
    variable r2241 : std_logic_vector(0 to 0) := (others => '0');
    variable r2240 : std_logic_vector(0 to 0) := (others => '0');
    variable r2239 : std_logic_vector(0 to 0) := (others => '0');
    variable r2238 : std_logic_vector(0 to 0) := (others => '0');
    variable r2237 : std_logic_vector(0 to 0) := (others => '0');
    variable r2236 : std_logic_vector(0 to 0) := (others => '0');
    variable r2235 : std_logic_vector(0 to 0) := (others => '0');
    variable r2234 : std_logic_vector(0 to 0) := (others => '0');
    variable r2233 : std_logic_vector(0 to 0) := (others => '0');
    variable r2232 : std_logic_vector(0 to 0) := (others => '0');
    variable r2231 : std_logic_vector(0 to 0) := (others => '0');
    variable r2230 : std_logic_vector(0 to 0) := (others => '0');
    variable r2229 : std_logic_vector(0 to 0) := (others => '0');
    variable r2228 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r2229 := "1";
    null;
    r2230 := (r2229);
    r2231 := "1";
    null;
    r2232 := (r2231);
    r2233 := "0";
    null;
    r2234 := (r2233);
    r2235 := "1";
    null;
    r2236 := (r2235);
    r2237 := "1";
    null;
    r2238 := (r2237);
    r2239 := "0";
    null;
    r2240 := (r2239);
    r2241 := "0";
    null;
    r2242 := (r2241);
    r2243 := "0";
    null;
    r2244 := (r2243);
    r2245 := "0";
    null;
    r2246 := (r2245);
    r2247 := "0";
    null;
    r2248 := (r2247);
    r2249 := "0";
    null;
    r2250 := (r2249);
    r2251 := "0";
    null;
    r2252 := (r2251);
    r2253 := "0";
    null;
    r2254 := (r2253);
    r2255 := "1";
    null;
    r2256 := (r2255);
    r2257 := "1";
    null;
    r2258 := (r2257);
    r2259 := "1";
    null;
    r2260 := (r2259);
    r2261 := "1";
    null;
    r2262 := (r2261);
    r2263 := "0";
    null;
    r2264 := (r2263);
    r2265 := "1";
    null;
    r2266 := (r2265);
    r2267 := "0";
    null;
    r2268 := (r2267);
    r2269 := "1";
    null;
    r2270 := (r2269);
    r2271 := "0";
    null;
    r2272 := (r2271);
    r2273 := "1";
    null;
    r2274 := (r2273);
    r2275 := "0";
    null;
    r2276 := (r2275);
    r2277 := "1";
    null;
    r2278 := (r2277);
    r2279 := "0";
    null;
    r2280 := (r2279);
    r2281 := "0";
    null;
    r2282 := (r2281);
    r2283 := "1";
    null;
    r2284 := (r2283);
    r2285 := "1";
    null;
    r2286 := (r2285);
    r2287 := "0";
    null;
    r2288 := (r2287);
    r2289 := "0";
    null;
    r2290 := (r2289);
    r2291 := "0";
    null;
    r2292 := (r2291);
    r2228 := (r2230 & r2232 & r2234 & r2236 & r2238 & r2240 & r2242 & r2244 & r2246 & r2248 & r2250 & r2252 & r2254 & r2256 & r2258 & r2260 & r2262 & r2264 & r2266 & r2268 & r2270 & r2272 & r2274 & r2276 & r2278 & r2280 & r2282 & r2284 & r2286 & r2288 & r2290 & r2292);
    return r2228;
  end rewire_MetaprogrammingRW.wd807aa98_2227;
  function rewire_MetaprogrammingRW.wab1c5ed5_2158 return std_logic_vector
  is
    variable r2223 : std_logic_vector(0 to 0) := (others => '0');
    variable r2222 : std_logic_vector(0 to 0) := (others => '0');
    variable r2221 : std_logic_vector(0 to 0) := (others => '0');
    variable r2220 : std_logic_vector(0 to 0) := (others => '0');
    variable r2219 : std_logic_vector(0 to 0) := (others => '0');
    variable r2218 : std_logic_vector(0 to 0) := (others => '0');
    variable r2217 : std_logic_vector(0 to 0) := (others => '0');
    variable r2216 : std_logic_vector(0 to 0) := (others => '0');
    variable r2215 : std_logic_vector(0 to 0) := (others => '0');
    variable r2214 : std_logic_vector(0 to 0) := (others => '0');
    variable r2213 : std_logic_vector(0 to 0) := (others => '0');
    variable r2212 : std_logic_vector(0 to 0) := (others => '0');
    variable r2211 : std_logic_vector(0 to 0) := (others => '0');
    variable r2210 : std_logic_vector(0 to 0) := (others => '0');
    variable r2209 : std_logic_vector(0 to 0) := (others => '0');
    variable r2208 : std_logic_vector(0 to 0) := (others => '0');
    variable r2207 : std_logic_vector(0 to 0) := (others => '0');
    variable r2206 : std_logic_vector(0 to 0) := (others => '0');
    variable r2205 : std_logic_vector(0 to 0) := (others => '0');
    variable r2204 : std_logic_vector(0 to 0) := (others => '0');
    variable r2203 : std_logic_vector(0 to 0) := (others => '0');
    variable r2202 : std_logic_vector(0 to 0) := (others => '0');
    variable r2201 : std_logic_vector(0 to 0) := (others => '0');
    variable r2200 : std_logic_vector(0 to 0) := (others => '0');
    variable r2199 : std_logic_vector(0 to 0) := (others => '0');
    variable r2198 : std_logic_vector(0 to 0) := (others => '0');
    variable r2197 : std_logic_vector(0 to 0) := (others => '0');
    variable r2196 : std_logic_vector(0 to 0) := (others => '0');
    variable r2195 : std_logic_vector(0 to 0) := (others => '0');
    variable r2194 : std_logic_vector(0 to 0) := (others => '0');
    variable r2193 : std_logic_vector(0 to 0) := (others => '0');
    variable r2192 : std_logic_vector(0 to 0) := (others => '0');
    variable r2191 : std_logic_vector(0 to 0) := (others => '0');
    variable r2190 : std_logic_vector(0 to 0) := (others => '0');
    variable r2189 : std_logic_vector(0 to 0) := (others => '0');
    variable r2188 : std_logic_vector(0 to 0) := (others => '0');
    variable r2187 : std_logic_vector(0 to 0) := (others => '0');
    variable r2186 : std_logic_vector(0 to 0) := (others => '0');
    variable r2185 : std_logic_vector(0 to 0) := (others => '0');
    variable r2184 : std_logic_vector(0 to 0) := (others => '0');
    variable r2183 : std_logic_vector(0 to 0) := (others => '0');
    variable r2182 : std_logic_vector(0 to 0) := (others => '0');
    variable r2181 : std_logic_vector(0 to 0) := (others => '0');
    variable r2180 : std_logic_vector(0 to 0) := (others => '0');
    variable r2179 : std_logic_vector(0 to 0) := (others => '0');
    variable r2178 : std_logic_vector(0 to 0) := (others => '0');
    variable r2177 : std_logic_vector(0 to 0) := (others => '0');
    variable r2176 : std_logic_vector(0 to 0) := (others => '0');
    variable r2175 : std_logic_vector(0 to 0) := (others => '0');
    variable r2174 : std_logic_vector(0 to 0) := (others => '0');
    variable r2173 : std_logic_vector(0 to 0) := (others => '0');
    variable r2172 : std_logic_vector(0 to 0) := (others => '0');
    variable r2171 : std_logic_vector(0 to 0) := (others => '0');
    variable r2170 : std_logic_vector(0 to 0) := (others => '0');
    variable r2169 : std_logic_vector(0 to 0) := (others => '0');
    variable r2168 : std_logic_vector(0 to 0) := (others => '0');
    variable r2167 : std_logic_vector(0 to 0) := (others => '0');
    variable r2166 : std_logic_vector(0 to 0) := (others => '0');
    variable r2165 : std_logic_vector(0 to 0) := (others => '0');
    variable r2164 : std_logic_vector(0 to 0) := (others => '0');
    variable r2163 : std_logic_vector(0 to 0) := (others => '0');
    variable r2162 : std_logic_vector(0 to 0) := (others => '0');
    variable r2161 : std_logic_vector(0 to 0) := (others => '0');
    variable r2160 : std_logic_vector(0 to 0) := (others => '0');
    variable r2159 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r2160 := "1";
    null;
    r2161 := (r2160);
    r2162 := "0";
    null;
    r2163 := (r2162);
    r2164 := "1";
    null;
    r2165 := (r2164);
    r2166 := "0";
    null;
    r2167 := (r2166);
    r2168 := "1";
    null;
    r2169 := (r2168);
    r2170 := "0";
    null;
    r2171 := (r2170);
    r2172 := "1";
    null;
    r2173 := (r2172);
    r2174 := "1";
    null;
    r2175 := (r2174);
    r2176 := "0";
    null;
    r2177 := (r2176);
    r2178 := "0";
    null;
    r2179 := (r2178);
    r2180 := "0";
    null;
    r2181 := (r2180);
    r2182 := "1";
    null;
    r2183 := (r2182);
    r2184 := "1";
    null;
    r2185 := (r2184);
    r2186 := "1";
    null;
    r2187 := (r2186);
    r2188 := "0";
    null;
    r2189 := (r2188);
    r2190 := "0";
    null;
    r2191 := (r2190);
    r2192 := "0";
    null;
    r2193 := (r2192);
    r2194 := "1";
    null;
    r2195 := (r2194);
    r2196 := "0";
    null;
    r2197 := (r2196);
    r2198 := "1";
    null;
    r2199 := (r2198);
    r2200 := "1";
    null;
    r2201 := (r2200);
    r2202 := "1";
    null;
    r2203 := (r2202);
    r2204 := "1";
    null;
    r2205 := (r2204);
    r2206 := "0";
    null;
    r2207 := (r2206);
    r2208 := "1";
    null;
    r2209 := (r2208);
    r2210 := "1";
    null;
    r2211 := (r2210);
    r2212 := "0";
    null;
    r2213 := (r2212);
    r2214 := "1";
    null;
    r2215 := (r2214);
    r2216 := "0";
    null;
    r2217 := (r2216);
    r2218 := "1";
    null;
    r2219 := (r2218);
    r2220 := "0";
    null;
    r2221 := (r2220);
    r2222 := "1";
    null;
    r2223 := (r2222);
    r2159 := (r2161 & r2163 & r2165 & r2167 & r2169 & r2171 & r2173 & r2175 & r2177 & r2179 & r2181 & r2183 & r2185 & r2187 & r2189 & r2191 & r2193 & r2195 & r2197 & r2199 & r2201 & r2203 & r2205 & r2207 & r2209 & r2211 & r2213 & r2215 & r2217 & r2219 & r2221 & r2223);
    return r2159;
  end rewire_MetaprogrammingRW.wab1c5ed5_2158;
  function rewire_MetaprogrammingRW.w923f82a4_2089 return std_logic_vector
  is
    variable r2154 : std_logic_vector(0 to 0) := (others => '0');
    variable r2153 : std_logic_vector(0 to 0) := (others => '0');
    variable r2152 : std_logic_vector(0 to 0) := (others => '0');
    variable r2151 : std_logic_vector(0 to 0) := (others => '0');
    variable r2150 : std_logic_vector(0 to 0) := (others => '0');
    variable r2149 : std_logic_vector(0 to 0) := (others => '0');
    variable r2148 : std_logic_vector(0 to 0) := (others => '0');
    variable r2147 : std_logic_vector(0 to 0) := (others => '0');
    variable r2146 : std_logic_vector(0 to 0) := (others => '0');
    variable r2145 : std_logic_vector(0 to 0) := (others => '0');
    variable r2144 : std_logic_vector(0 to 0) := (others => '0');
    variable r2143 : std_logic_vector(0 to 0) := (others => '0');
    variable r2142 : std_logic_vector(0 to 0) := (others => '0');
    variable r2141 : std_logic_vector(0 to 0) := (others => '0');
    variable r2140 : std_logic_vector(0 to 0) := (others => '0');
    variable r2139 : std_logic_vector(0 to 0) := (others => '0');
    variable r2138 : std_logic_vector(0 to 0) := (others => '0');
    variable r2137 : std_logic_vector(0 to 0) := (others => '0');
    variable r2136 : std_logic_vector(0 to 0) := (others => '0');
    variable r2135 : std_logic_vector(0 to 0) := (others => '0');
    variable r2134 : std_logic_vector(0 to 0) := (others => '0');
    variable r2133 : std_logic_vector(0 to 0) := (others => '0');
    variable r2132 : std_logic_vector(0 to 0) := (others => '0');
    variable r2131 : std_logic_vector(0 to 0) := (others => '0');
    variable r2130 : std_logic_vector(0 to 0) := (others => '0');
    variable r2129 : std_logic_vector(0 to 0) := (others => '0');
    variable r2128 : std_logic_vector(0 to 0) := (others => '0');
    variable r2127 : std_logic_vector(0 to 0) := (others => '0');
    variable r2126 : std_logic_vector(0 to 0) := (others => '0');
    variable r2125 : std_logic_vector(0 to 0) := (others => '0');
    variable r2124 : std_logic_vector(0 to 0) := (others => '0');
    variable r2123 : std_logic_vector(0 to 0) := (others => '0');
    variable r2122 : std_logic_vector(0 to 0) := (others => '0');
    variable r2121 : std_logic_vector(0 to 0) := (others => '0');
    variable r2120 : std_logic_vector(0 to 0) := (others => '0');
    variable r2119 : std_logic_vector(0 to 0) := (others => '0');
    variable r2118 : std_logic_vector(0 to 0) := (others => '0');
    variable r2117 : std_logic_vector(0 to 0) := (others => '0');
    variable r2116 : std_logic_vector(0 to 0) := (others => '0');
    variable r2115 : std_logic_vector(0 to 0) := (others => '0');
    variable r2114 : std_logic_vector(0 to 0) := (others => '0');
    variable r2113 : std_logic_vector(0 to 0) := (others => '0');
    variable r2112 : std_logic_vector(0 to 0) := (others => '0');
    variable r2111 : std_logic_vector(0 to 0) := (others => '0');
    variable r2110 : std_logic_vector(0 to 0) := (others => '0');
    variable r2109 : std_logic_vector(0 to 0) := (others => '0');
    variable r2108 : std_logic_vector(0 to 0) := (others => '0');
    variable r2107 : std_logic_vector(0 to 0) := (others => '0');
    variable r2106 : std_logic_vector(0 to 0) := (others => '0');
    variable r2105 : std_logic_vector(0 to 0) := (others => '0');
    variable r2104 : std_logic_vector(0 to 0) := (others => '0');
    variable r2103 : std_logic_vector(0 to 0) := (others => '0');
    variable r2102 : std_logic_vector(0 to 0) := (others => '0');
    variable r2101 : std_logic_vector(0 to 0) := (others => '0');
    variable r2100 : std_logic_vector(0 to 0) := (others => '0');
    variable r2099 : std_logic_vector(0 to 0) := (others => '0');
    variable r2098 : std_logic_vector(0 to 0) := (others => '0');
    variable r2097 : std_logic_vector(0 to 0) := (others => '0');
    variable r2096 : std_logic_vector(0 to 0) := (others => '0');
    variable r2095 : std_logic_vector(0 to 0) := (others => '0');
    variable r2094 : std_logic_vector(0 to 0) := (others => '0');
    variable r2093 : std_logic_vector(0 to 0) := (others => '0');
    variable r2092 : std_logic_vector(0 to 0) := (others => '0');
    variable r2091 : std_logic_vector(0 to 0) := (others => '0');
    variable r2090 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r2091 := "1";
    null;
    r2092 := (r2091);
    r2093 := "0";
    null;
    r2094 := (r2093);
    r2095 := "0";
    null;
    r2096 := (r2095);
    r2097 := "1";
    null;
    r2098 := (r2097);
    r2099 := "0";
    null;
    r2100 := (r2099);
    r2101 := "0";
    null;
    r2102 := (r2101);
    r2103 := "1";
    null;
    r2104 := (r2103);
    r2105 := "0";
    null;
    r2106 := (r2105);
    r2107 := "0";
    null;
    r2108 := (r2107);
    r2109 := "0";
    null;
    r2110 := (r2109);
    r2111 := "1";
    null;
    r2112 := (r2111);
    r2113 := "1";
    null;
    r2114 := (r2113);
    r2115 := "1";
    null;
    r2116 := (r2115);
    r2117 := "1";
    null;
    r2118 := (r2117);
    r2119 := "1";
    null;
    r2120 := (r2119);
    r2121 := "1";
    null;
    r2122 := (r2121);
    r2123 := "1";
    null;
    r2124 := (r2123);
    r2125 := "0";
    null;
    r2126 := (r2125);
    r2127 := "0";
    null;
    r2128 := (r2127);
    r2129 := "0";
    null;
    r2130 := (r2129);
    r2131 := "0";
    null;
    r2132 := (r2131);
    r2133 := "0";
    null;
    r2134 := (r2133);
    r2135 := "1";
    null;
    r2136 := (r2135);
    r2137 := "0";
    null;
    r2138 := (r2137);
    r2139 := "1";
    null;
    r2140 := (r2139);
    r2141 := "0";
    null;
    r2142 := (r2141);
    r2143 := "1";
    null;
    r2144 := (r2143);
    r2145 := "0";
    null;
    r2146 := (r2145);
    r2147 := "0";
    null;
    r2148 := (r2147);
    r2149 := "1";
    null;
    r2150 := (r2149);
    r2151 := "0";
    null;
    r2152 := (r2151);
    r2153 := "0";
    null;
    r2154 := (r2153);
    r2090 := (r2092 & r2094 & r2096 & r2098 & r2100 & r2102 & r2104 & r2106 & r2108 & r2110 & r2112 & r2114 & r2116 & r2118 & r2120 & r2122 & r2124 & r2126 & r2128 & r2130 & r2132 & r2134 & r2136 & r2138 & r2140 & r2142 & r2144 & r2146 & r2148 & r2150 & r2152 & r2154);
    return r2090;
  end rewire_MetaprogrammingRW.w923f82a4_2089;
  function rewire_MetaprogrammingRW.w59f111f1_2020 return std_logic_vector
  is
    variable r2085 : std_logic_vector(0 to 0) := (others => '0');
    variable r2084 : std_logic_vector(0 to 0) := (others => '0');
    variable r2083 : std_logic_vector(0 to 0) := (others => '0');
    variable r2082 : std_logic_vector(0 to 0) := (others => '0');
    variable r2081 : std_logic_vector(0 to 0) := (others => '0');
    variable r2080 : std_logic_vector(0 to 0) := (others => '0');
    variable r2079 : std_logic_vector(0 to 0) := (others => '0');
    variable r2078 : std_logic_vector(0 to 0) := (others => '0');
    variable r2077 : std_logic_vector(0 to 0) := (others => '0');
    variable r2076 : std_logic_vector(0 to 0) := (others => '0');
    variable r2075 : std_logic_vector(0 to 0) := (others => '0');
    variable r2074 : std_logic_vector(0 to 0) := (others => '0');
    variable r2073 : std_logic_vector(0 to 0) := (others => '0');
    variable r2072 : std_logic_vector(0 to 0) := (others => '0');
    variable r2071 : std_logic_vector(0 to 0) := (others => '0');
    variable r2070 : std_logic_vector(0 to 0) := (others => '0');
    variable r2069 : std_logic_vector(0 to 0) := (others => '0');
    variable r2068 : std_logic_vector(0 to 0) := (others => '0');
    variable r2067 : std_logic_vector(0 to 0) := (others => '0');
    variable r2066 : std_logic_vector(0 to 0) := (others => '0');
    variable r2065 : std_logic_vector(0 to 0) := (others => '0');
    variable r2064 : std_logic_vector(0 to 0) := (others => '0');
    variable r2063 : std_logic_vector(0 to 0) := (others => '0');
    variable r2062 : std_logic_vector(0 to 0) := (others => '0');
    variable r2061 : std_logic_vector(0 to 0) := (others => '0');
    variable r2060 : std_logic_vector(0 to 0) := (others => '0');
    variable r2059 : std_logic_vector(0 to 0) := (others => '0');
    variable r2058 : std_logic_vector(0 to 0) := (others => '0');
    variable r2057 : std_logic_vector(0 to 0) := (others => '0');
    variable r2056 : std_logic_vector(0 to 0) := (others => '0');
    variable r2055 : std_logic_vector(0 to 0) := (others => '0');
    variable r2054 : std_logic_vector(0 to 0) := (others => '0');
    variable r2053 : std_logic_vector(0 to 0) := (others => '0');
    variable r2052 : std_logic_vector(0 to 0) := (others => '0');
    variable r2051 : std_logic_vector(0 to 0) := (others => '0');
    variable r2050 : std_logic_vector(0 to 0) := (others => '0');
    variable r2049 : std_logic_vector(0 to 0) := (others => '0');
    variable r2048 : std_logic_vector(0 to 0) := (others => '0');
    variable r2047 : std_logic_vector(0 to 0) := (others => '0');
    variable r2046 : std_logic_vector(0 to 0) := (others => '0');
    variable r2045 : std_logic_vector(0 to 0) := (others => '0');
    variable r2044 : std_logic_vector(0 to 0) := (others => '0');
    variable r2043 : std_logic_vector(0 to 0) := (others => '0');
    variable r2042 : std_logic_vector(0 to 0) := (others => '0');
    variable r2041 : std_logic_vector(0 to 0) := (others => '0');
    variable r2040 : std_logic_vector(0 to 0) := (others => '0');
    variable r2039 : std_logic_vector(0 to 0) := (others => '0');
    variable r2038 : std_logic_vector(0 to 0) := (others => '0');
    variable r2037 : std_logic_vector(0 to 0) := (others => '0');
    variable r2036 : std_logic_vector(0 to 0) := (others => '0');
    variable r2035 : std_logic_vector(0 to 0) := (others => '0');
    variable r2034 : std_logic_vector(0 to 0) := (others => '0');
    variable r2033 : std_logic_vector(0 to 0) := (others => '0');
    variable r2032 : std_logic_vector(0 to 0) := (others => '0');
    variable r2031 : std_logic_vector(0 to 0) := (others => '0');
    variable r2030 : std_logic_vector(0 to 0) := (others => '0');
    variable r2029 : std_logic_vector(0 to 0) := (others => '0');
    variable r2028 : std_logic_vector(0 to 0) := (others => '0');
    variable r2027 : std_logic_vector(0 to 0) := (others => '0');
    variable r2026 : std_logic_vector(0 to 0) := (others => '0');
    variable r2025 : std_logic_vector(0 to 0) := (others => '0');
    variable r2024 : std_logic_vector(0 to 0) := (others => '0');
    variable r2023 : std_logic_vector(0 to 0) := (others => '0');
    variable r2022 : std_logic_vector(0 to 0) := (others => '0');
    variable r2021 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r2022 := "0";
    null;
    r2023 := (r2022);
    r2024 := "1";
    null;
    r2025 := (r2024);
    r2026 := "0";
    null;
    r2027 := (r2026);
    r2028 := "1";
    null;
    r2029 := (r2028);
    r2030 := "1";
    null;
    r2031 := (r2030);
    r2032 := "0";
    null;
    r2033 := (r2032);
    r2034 := "0";
    null;
    r2035 := (r2034);
    r2036 := "1";
    null;
    r2037 := (r2036);
    r2038 := "1";
    null;
    r2039 := (r2038);
    r2040 := "1";
    null;
    r2041 := (r2040);
    r2042 := "1";
    null;
    r2043 := (r2042);
    r2044 := "1";
    null;
    r2045 := (r2044);
    r2046 := "0";
    null;
    r2047 := (r2046);
    r2048 := "0";
    null;
    r2049 := (r2048);
    r2050 := "0";
    null;
    r2051 := (r2050);
    r2052 := "1";
    null;
    r2053 := (r2052);
    r2054 := "0";
    null;
    r2055 := (r2054);
    r2056 := "0";
    null;
    r2057 := (r2056);
    r2058 := "0";
    null;
    r2059 := (r2058);
    r2060 := "1";
    null;
    r2061 := (r2060);
    r2062 := "0";
    null;
    r2063 := (r2062);
    r2064 := "0";
    null;
    r2065 := (r2064);
    r2066 := "0";
    null;
    r2067 := (r2066);
    r2068 := "1";
    null;
    r2069 := (r2068);
    r2070 := "1";
    null;
    r2071 := (r2070);
    r2072 := "1";
    null;
    r2073 := (r2072);
    r2074 := "1";
    null;
    r2075 := (r2074);
    r2076 := "1";
    null;
    r2077 := (r2076);
    r2078 := "0";
    null;
    r2079 := (r2078);
    r2080 := "0";
    null;
    r2081 := (r2080);
    r2082 := "0";
    null;
    r2083 := (r2082);
    r2084 := "1";
    null;
    r2085 := (r2084);
    r2021 := (r2023 & r2025 & r2027 & r2029 & r2031 & r2033 & r2035 & r2037 & r2039 & r2041 & r2043 & r2045 & r2047 & r2049 & r2051 & r2053 & r2055 & r2057 & r2059 & r2061 & r2063 & r2065 & r2067 & r2069 & r2071 & r2073 & r2075 & r2077 & r2079 & r2081 & r2083 & r2085);
    return r2021;
  end rewire_MetaprogrammingRW.w59f111f1_2020;
  function rewire_MetaprogrammingRW.w3956c25b_1951 return std_logic_vector
  is
    variable r2016 : std_logic_vector(0 to 0) := (others => '0');
    variable r2015 : std_logic_vector(0 to 0) := (others => '0');
    variable r2014 : std_logic_vector(0 to 0) := (others => '0');
    variable r2013 : std_logic_vector(0 to 0) := (others => '0');
    variable r2012 : std_logic_vector(0 to 0) := (others => '0');
    variable r2011 : std_logic_vector(0 to 0) := (others => '0');
    variable r2010 : std_logic_vector(0 to 0) := (others => '0');
    variable r2009 : std_logic_vector(0 to 0) := (others => '0');
    variable r2008 : std_logic_vector(0 to 0) := (others => '0');
    variable r2007 : std_logic_vector(0 to 0) := (others => '0');
    variable r2006 : std_logic_vector(0 to 0) := (others => '0');
    variable r2005 : std_logic_vector(0 to 0) := (others => '0');
    variable r2004 : std_logic_vector(0 to 0) := (others => '0');
    variable r2003 : std_logic_vector(0 to 0) := (others => '0');
    variable r2002 : std_logic_vector(0 to 0) := (others => '0');
    variable r2001 : std_logic_vector(0 to 0) := (others => '0');
    variable r2000 : std_logic_vector(0 to 0) := (others => '0');
    variable r1999 : std_logic_vector(0 to 0) := (others => '0');
    variable r1998 : std_logic_vector(0 to 0) := (others => '0');
    variable r1997 : std_logic_vector(0 to 0) := (others => '0');
    variable r1996 : std_logic_vector(0 to 0) := (others => '0');
    variable r1995 : std_logic_vector(0 to 0) := (others => '0');
    variable r1994 : std_logic_vector(0 to 0) := (others => '0');
    variable r1993 : std_logic_vector(0 to 0) := (others => '0');
    variable r1992 : std_logic_vector(0 to 0) := (others => '0');
    variable r1991 : std_logic_vector(0 to 0) := (others => '0');
    variable r1990 : std_logic_vector(0 to 0) := (others => '0');
    variable r1989 : std_logic_vector(0 to 0) := (others => '0');
    variable r1988 : std_logic_vector(0 to 0) := (others => '0');
    variable r1987 : std_logic_vector(0 to 0) := (others => '0');
    variable r1986 : std_logic_vector(0 to 0) := (others => '0');
    variable r1985 : std_logic_vector(0 to 0) := (others => '0');
    variable r1984 : std_logic_vector(0 to 0) := (others => '0');
    variable r1983 : std_logic_vector(0 to 0) := (others => '0');
    variable r1982 : std_logic_vector(0 to 0) := (others => '0');
    variable r1981 : std_logic_vector(0 to 0) := (others => '0');
    variable r1980 : std_logic_vector(0 to 0) := (others => '0');
    variable r1979 : std_logic_vector(0 to 0) := (others => '0');
    variable r1978 : std_logic_vector(0 to 0) := (others => '0');
    variable r1977 : std_logic_vector(0 to 0) := (others => '0');
    variable r1976 : std_logic_vector(0 to 0) := (others => '0');
    variable r1975 : std_logic_vector(0 to 0) := (others => '0');
    variable r1974 : std_logic_vector(0 to 0) := (others => '0');
    variable r1973 : std_logic_vector(0 to 0) := (others => '0');
    variable r1972 : std_logic_vector(0 to 0) := (others => '0');
    variable r1971 : std_logic_vector(0 to 0) := (others => '0');
    variable r1970 : std_logic_vector(0 to 0) := (others => '0');
    variable r1969 : std_logic_vector(0 to 0) := (others => '0');
    variable r1968 : std_logic_vector(0 to 0) := (others => '0');
    variable r1967 : std_logic_vector(0 to 0) := (others => '0');
    variable r1966 : std_logic_vector(0 to 0) := (others => '0');
    variable r1965 : std_logic_vector(0 to 0) := (others => '0');
    variable r1964 : std_logic_vector(0 to 0) := (others => '0');
    variable r1963 : std_logic_vector(0 to 0) := (others => '0');
    variable r1962 : std_logic_vector(0 to 0) := (others => '0');
    variable r1961 : std_logic_vector(0 to 0) := (others => '0');
    variable r1960 : std_logic_vector(0 to 0) := (others => '0');
    variable r1959 : std_logic_vector(0 to 0) := (others => '0');
    variable r1958 : std_logic_vector(0 to 0) := (others => '0');
    variable r1957 : std_logic_vector(0 to 0) := (others => '0');
    variable r1956 : std_logic_vector(0 to 0) := (others => '0');
    variable r1955 : std_logic_vector(0 to 0) := (others => '0');
    variable r1954 : std_logic_vector(0 to 0) := (others => '0');
    variable r1953 : std_logic_vector(0 to 0) := (others => '0');
    variable r1952 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r1953 := "0";
    null;
    r1954 := (r1953);
    r1955 := "0";
    null;
    r1956 := (r1955);
    r1957 := "1";
    null;
    r1958 := (r1957);
    r1959 := "1";
    null;
    r1960 := (r1959);
    r1961 := "1";
    null;
    r1962 := (r1961);
    r1963 := "0";
    null;
    r1964 := (r1963);
    r1965 := "0";
    null;
    r1966 := (r1965);
    r1967 := "1";
    null;
    r1968 := (r1967);
    r1969 := "0";
    null;
    r1970 := (r1969);
    r1971 := "1";
    null;
    r1972 := (r1971);
    r1973 := "0";
    null;
    r1974 := (r1973);
    r1975 := "1";
    null;
    r1976 := (r1975);
    r1977 := "0";
    null;
    r1978 := (r1977);
    r1979 := "1";
    null;
    r1980 := (r1979);
    r1981 := "1";
    null;
    r1982 := (r1981);
    r1983 := "0";
    null;
    r1984 := (r1983);
    r1985 := "1";
    null;
    r1986 := (r1985);
    r1987 := "1";
    null;
    r1988 := (r1987);
    r1989 := "0";
    null;
    r1990 := (r1989);
    r1991 := "0";
    null;
    r1992 := (r1991);
    r1993 := "0";
    null;
    r1994 := (r1993);
    r1995 := "0";
    null;
    r1996 := (r1995);
    r1997 := "1";
    null;
    r1998 := (r1997);
    r1999 := "0";
    null;
    r2000 := (r1999);
    r2001 := "0";
    null;
    r2002 := (r2001);
    r2003 := "1";
    null;
    r2004 := (r2003);
    r2005 := "0";
    null;
    r2006 := (r2005);
    r2007 := "1";
    null;
    r2008 := (r2007);
    r2009 := "1";
    null;
    r2010 := (r2009);
    r2011 := "0";
    null;
    r2012 := (r2011);
    r2013 := "1";
    null;
    r2014 := (r2013);
    r2015 := "1";
    null;
    r2016 := (r2015);
    r1952 := (r1954 & r1956 & r1958 & r1960 & r1962 & r1964 & r1966 & r1968 & r1970 & r1972 & r1974 & r1976 & r1978 & r1980 & r1982 & r1984 & r1986 & r1988 & r1990 & r1992 & r1994 & r1996 & r1998 & r2000 & r2002 & r2004 & r2006 & r2008 & r2010 & r2012 & r2014 & r2016);
    return r1952;
  end rewire_MetaprogrammingRW.w3956c25b_1951;
  function rewire_MetaprogrammingRW.we9b5dba5_1882 return std_logic_vector
  is
    variable r1947 : std_logic_vector(0 to 0) := (others => '0');
    variable r1946 : std_logic_vector(0 to 0) := (others => '0');
    variable r1945 : std_logic_vector(0 to 0) := (others => '0');
    variable r1944 : std_logic_vector(0 to 0) := (others => '0');
    variable r1943 : std_logic_vector(0 to 0) := (others => '0');
    variable r1942 : std_logic_vector(0 to 0) := (others => '0');
    variable r1941 : std_logic_vector(0 to 0) := (others => '0');
    variable r1940 : std_logic_vector(0 to 0) := (others => '0');
    variable r1939 : std_logic_vector(0 to 0) := (others => '0');
    variable r1938 : std_logic_vector(0 to 0) := (others => '0');
    variable r1937 : std_logic_vector(0 to 0) := (others => '0');
    variable r1936 : std_logic_vector(0 to 0) := (others => '0');
    variable r1935 : std_logic_vector(0 to 0) := (others => '0');
    variable r1934 : std_logic_vector(0 to 0) := (others => '0');
    variable r1933 : std_logic_vector(0 to 0) := (others => '0');
    variable r1932 : std_logic_vector(0 to 0) := (others => '0');
    variable r1931 : std_logic_vector(0 to 0) := (others => '0');
    variable r1930 : std_logic_vector(0 to 0) := (others => '0');
    variable r1929 : std_logic_vector(0 to 0) := (others => '0');
    variable r1928 : std_logic_vector(0 to 0) := (others => '0');
    variable r1927 : std_logic_vector(0 to 0) := (others => '0');
    variable r1926 : std_logic_vector(0 to 0) := (others => '0');
    variable r1925 : std_logic_vector(0 to 0) := (others => '0');
    variable r1924 : std_logic_vector(0 to 0) := (others => '0');
    variable r1923 : std_logic_vector(0 to 0) := (others => '0');
    variable r1922 : std_logic_vector(0 to 0) := (others => '0');
    variable r1921 : std_logic_vector(0 to 0) := (others => '0');
    variable r1920 : std_logic_vector(0 to 0) := (others => '0');
    variable r1919 : std_logic_vector(0 to 0) := (others => '0');
    variable r1918 : std_logic_vector(0 to 0) := (others => '0');
    variable r1917 : std_logic_vector(0 to 0) := (others => '0');
    variable r1916 : std_logic_vector(0 to 0) := (others => '0');
    variable r1915 : std_logic_vector(0 to 0) := (others => '0');
    variable r1914 : std_logic_vector(0 to 0) := (others => '0');
    variable r1913 : std_logic_vector(0 to 0) := (others => '0');
    variable r1912 : std_logic_vector(0 to 0) := (others => '0');
    variable r1911 : std_logic_vector(0 to 0) := (others => '0');
    variable r1910 : std_logic_vector(0 to 0) := (others => '0');
    variable r1909 : std_logic_vector(0 to 0) := (others => '0');
    variable r1908 : std_logic_vector(0 to 0) := (others => '0');
    variable r1907 : std_logic_vector(0 to 0) := (others => '0');
    variable r1906 : std_logic_vector(0 to 0) := (others => '0');
    variable r1905 : std_logic_vector(0 to 0) := (others => '0');
    variable r1904 : std_logic_vector(0 to 0) := (others => '0');
    variable r1903 : std_logic_vector(0 to 0) := (others => '0');
    variable r1902 : std_logic_vector(0 to 0) := (others => '0');
    variable r1901 : std_logic_vector(0 to 0) := (others => '0');
    variable r1900 : std_logic_vector(0 to 0) := (others => '0');
    variable r1899 : std_logic_vector(0 to 0) := (others => '0');
    variable r1898 : std_logic_vector(0 to 0) := (others => '0');
    variable r1897 : std_logic_vector(0 to 0) := (others => '0');
    variable r1896 : std_logic_vector(0 to 0) := (others => '0');
    variable r1895 : std_logic_vector(0 to 0) := (others => '0');
    variable r1894 : std_logic_vector(0 to 0) := (others => '0');
    variable r1893 : std_logic_vector(0 to 0) := (others => '0');
    variable r1892 : std_logic_vector(0 to 0) := (others => '0');
    variable r1891 : std_logic_vector(0 to 0) := (others => '0');
    variable r1890 : std_logic_vector(0 to 0) := (others => '0');
    variable r1889 : std_logic_vector(0 to 0) := (others => '0');
    variable r1888 : std_logic_vector(0 to 0) := (others => '0');
    variable r1887 : std_logic_vector(0 to 0) := (others => '0');
    variable r1886 : std_logic_vector(0 to 0) := (others => '0');
    variable r1885 : std_logic_vector(0 to 0) := (others => '0');
    variable r1884 : std_logic_vector(0 to 0) := (others => '0');
    variable r1883 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r1884 := "1";
    null;
    r1885 := (r1884);
    r1886 := "1";
    null;
    r1887 := (r1886);
    r1888 := "1";
    null;
    r1889 := (r1888);
    r1890 := "0";
    null;
    r1891 := (r1890);
    r1892 := "1";
    null;
    r1893 := (r1892);
    r1894 := "0";
    null;
    r1895 := (r1894);
    r1896 := "0";
    null;
    r1897 := (r1896);
    r1898 := "1";
    null;
    r1899 := (r1898);
    r1900 := "1";
    null;
    r1901 := (r1900);
    r1902 := "0";
    null;
    r1903 := (r1902);
    r1904 := "1";
    null;
    r1905 := (r1904);
    r1906 := "1";
    null;
    r1907 := (r1906);
    r1908 := "0";
    null;
    r1909 := (r1908);
    r1910 := "1";
    null;
    r1911 := (r1910);
    r1912 := "0";
    null;
    r1913 := (r1912);
    r1914 := "1";
    null;
    r1915 := (r1914);
    r1916 := "1";
    null;
    r1917 := (r1916);
    r1918 := "1";
    null;
    r1919 := (r1918);
    r1920 := "0";
    null;
    r1921 := (r1920);
    r1922 := "1";
    null;
    r1923 := (r1922);
    r1924 := "1";
    null;
    r1925 := (r1924);
    r1926 := "0";
    null;
    r1927 := (r1926);
    r1928 := "1";
    null;
    r1929 := (r1928);
    r1930 := "1";
    null;
    r1931 := (r1930);
    r1932 := "1";
    null;
    r1933 := (r1932);
    r1934 := "0";
    null;
    r1935 := (r1934);
    r1936 := "1";
    null;
    r1937 := (r1936);
    r1938 := "0";
    null;
    r1939 := (r1938);
    r1940 := "0";
    null;
    r1941 := (r1940);
    r1942 := "1";
    null;
    r1943 := (r1942);
    r1944 := "0";
    null;
    r1945 := (r1944);
    r1946 := "1";
    null;
    r1947 := (r1946);
    r1883 := (r1885 & r1887 & r1889 & r1891 & r1893 & r1895 & r1897 & r1899 & r1901 & r1903 & r1905 & r1907 & r1909 & r1911 & r1913 & r1915 & r1917 & r1919 & r1921 & r1923 & r1925 & r1927 & r1929 & r1931 & r1933 & r1935 & r1937 & r1939 & r1941 & r1943 & r1945 & r1947);
    return r1883;
  end rewire_MetaprogrammingRW.we9b5dba5_1882;
  function rewire_MetaprogrammingRW.wb5c0fbcf_1813 return std_logic_vector
  is
    variable r1878 : std_logic_vector(0 to 0) := (others => '0');
    variable r1877 : std_logic_vector(0 to 0) := (others => '0');
    variable r1876 : std_logic_vector(0 to 0) := (others => '0');
    variable r1875 : std_logic_vector(0 to 0) := (others => '0');
    variable r1874 : std_logic_vector(0 to 0) := (others => '0');
    variable r1873 : std_logic_vector(0 to 0) := (others => '0');
    variable r1872 : std_logic_vector(0 to 0) := (others => '0');
    variable r1871 : std_logic_vector(0 to 0) := (others => '0');
    variable r1870 : std_logic_vector(0 to 0) := (others => '0');
    variable r1869 : std_logic_vector(0 to 0) := (others => '0');
    variable r1868 : std_logic_vector(0 to 0) := (others => '0');
    variable r1867 : std_logic_vector(0 to 0) := (others => '0');
    variable r1866 : std_logic_vector(0 to 0) := (others => '0');
    variable r1865 : std_logic_vector(0 to 0) := (others => '0');
    variable r1864 : std_logic_vector(0 to 0) := (others => '0');
    variable r1863 : std_logic_vector(0 to 0) := (others => '0');
    variable r1862 : std_logic_vector(0 to 0) := (others => '0');
    variable r1861 : std_logic_vector(0 to 0) := (others => '0');
    variable r1860 : std_logic_vector(0 to 0) := (others => '0');
    variable r1859 : std_logic_vector(0 to 0) := (others => '0');
    variable r1858 : std_logic_vector(0 to 0) := (others => '0');
    variable r1857 : std_logic_vector(0 to 0) := (others => '0');
    variable r1856 : std_logic_vector(0 to 0) := (others => '0');
    variable r1855 : std_logic_vector(0 to 0) := (others => '0');
    variable r1854 : std_logic_vector(0 to 0) := (others => '0');
    variable r1853 : std_logic_vector(0 to 0) := (others => '0');
    variable r1852 : std_logic_vector(0 to 0) := (others => '0');
    variable r1851 : std_logic_vector(0 to 0) := (others => '0');
    variable r1850 : std_logic_vector(0 to 0) := (others => '0');
    variable r1849 : std_logic_vector(0 to 0) := (others => '0');
    variable r1848 : std_logic_vector(0 to 0) := (others => '0');
    variable r1847 : std_logic_vector(0 to 0) := (others => '0');
    variable r1846 : std_logic_vector(0 to 0) := (others => '0');
    variable r1845 : std_logic_vector(0 to 0) := (others => '0');
    variable r1844 : std_logic_vector(0 to 0) := (others => '0');
    variable r1843 : std_logic_vector(0 to 0) := (others => '0');
    variable r1842 : std_logic_vector(0 to 0) := (others => '0');
    variable r1841 : std_logic_vector(0 to 0) := (others => '0');
    variable r1840 : std_logic_vector(0 to 0) := (others => '0');
    variable r1839 : std_logic_vector(0 to 0) := (others => '0');
    variable r1838 : std_logic_vector(0 to 0) := (others => '0');
    variable r1837 : std_logic_vector(0 to 0) := (others => '0');
    variable r1836 : std_logic_vector(0 to 0) := (others => '0');
    variable r1835 : std_logic_vector(0 to 0) := (others => '0');
    variable r1834 : std_logic_vector(0 to 0) := (others => '0');
    variable r1833 : std_logic_vector(0 to 0) := (others => '0');
    variable r1832 : std_logic_vector(0 to 0) := (others => '0');
    variable r1831 : std_logic_vector(0 to 0) := (others => '0');
    variable r1830 : std_logic_vector(0 to 0) := (others => '0');
    variable r1829 : std_logic_vector(0 to 0) := (others => '0');
    variable r1828 : std_logic_vector(0 to 0) := (others => '0');
    variable r1827 : std_logic_vector(0 to 0) := (others => '0');
    variable r1826 : std_logic_vector(0 to 0) := (others => '0');
    variable r1825 : std_logic_vector(0 to 0) := (others => '0');
    variable r1824 : std_logic_vector(0 to 0) := (others => '0');
    variable r1823 : std_logic_vector(0 to 0) := (others => '0');
    variable r1822 : std_logic_vector(0 to 0) := (others => '0');
    variable r1821 : std_logic_vector(0 to 0) := (others => '0');
    variable r1820 : std_logic_vector(0 to 0) := (others => '0');
    variable r1819 : std_logic_vector(0 to 0) := (others => '0');
    variable r1818 : std_logic_vector(0 to 0) := (others => '0');
    variable r1817 : std_logic_vector(0 to 0) := (others => '0');
    variable r1816 : std_logic_vector(0 to 0) := (others => '0');
    variable r1815 : std_logic_vector(0 to 0) := (others => '0');
    variable r1814 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r1815 := "1";
    null;
    r1816 := (r1815);
    r1817 := "0";
    null;
    r1818 := (r1817);
    r1819 := "1";
    null;
    r1820 := (r1819);
    r1821 := "1";
    null;
    r1822 := (r1821);
    r1823 := "0";
    null;
    r1824 := (r1823);
    r1825 := "1";
    null;
    r1826 := (r1825);
    r1827 := "0";
    null;
    r1828 := (r1827);
    r1829 := "1";
    null;
    r1830 := (r1829);
    r1831 := "1";
    null;
    r1832 := (r1831);
    r1833 := "1";
    null;
    r1834 := (r1833);
    r1835 := "0";
    null;
    r1836 := (r1835);
    r1837 := "0";
    null;
    r1838 := (r1837);
    r1839 := "0";
    null;
    r1840 := (r1839);
    r1841 := "0";
    null;
    r1842 := (r1841);
    r1843 := "0";
    null;
    r1844 := (r1843);
    r1845 := "0";
    null;
    r1846 := (r1845);
    r1847 := "1";
    null;
    r1848 := (r1847);
    r1849 := "1";
    null;
    r1850 := (r1849);
    r1851 := "1";
    null;
    r1852 := (r1851);
    r1853 := "1";
    null;
    r1854 := (r1853);
    r1855 := "1";
    null;
    r1856 := (r1855);
    r1857 := "0";
    null;
    r1858 := (r1857);
    r1859 := "1";
    null;
    r1860 := (r1859);
    r1861 := "1";
    null;
    r1862 := (r1861);
    r1863 := "1";
    null;
    r1864 := (r1863);
    r1865 := "1";
    null;
    r1866 := (r1865);
    r1867 := "0";
    null;
    r1868 := (r1867);
    r1869 := "0";
    null;
    r1870 := (r1869);
    r1871 := "1";
    null;
    r1872 := (r1871);
    r1873 := "1";
    null;
    r1874 := (r1873);
    r1875 := "1";
    null;
    r1876 := (r1875);
    r1877 := "1";
    null;
    r1878 := (r1877);
    r1814 := (r1816 & r1818 & r1820 & r1822 & r1824 & r1826 & r1828 & r1830 & r1832 & r1834 & r1836 & r1838 & r1840 & r1842 & r1844 & r1846 & r1848 & r1850 & r1852 & r1854 & r1856 & r1858 & r1860 & r1862 & r1864 & r1866 & r1868 & r1870 & r1872 & r1874 & r1876 & r1878);
    return r1814;
  end rewire_MetaprogrammingRW.wb5c0fbcf_1813;
  function rewire_MetaprogrammingRW.w71374491_1744 return std_logic_vector
  is
    variable r1809 : std_logic_vector(0 to 0) := (others => '0');
    variable r1808 : std_logic_vector(0 to 0) := (others => '0');
    variable r1807 : std_logic_vector(0 to 0) := (others => '0');
    variable r1806 : std_logic_vector(0 to 0) := (others => '0');
    variable r1805 : std_logic_vector(0 to 0) := (others => '0');
    variable r1804 : std_logic_vector(0 to 0) := (others => '0');
    variable r1803 : std_logic_vector(0 to 0) := (others => '0');
    variable r1802 : std_logic_vector(0 to 0) := (others => '0');
    variable r1801 : std_logic_vector(0 to 0) := (others => '0');
    variable r1800 : std_logic_vector(0 to 0) := (others => '0');
    variable r1799 : std_logic_vector(0 to 0) := (others => '0');
    variable r1798 : std_logic_vector(0 to 0) := (others => '0');
    variable r1797 : std_logic_vector(0 to 0) := (others => '0');
    variable r1796 : std_logic_vector(0 to 0) := (others => '0');
    variable r1795 : std_logic_vector(0 to 0) := (others => '0');
    variable r1794 : std_logic_vector(0 to 0) := (others => '0');
    variable r1793 : std_logic_vector(0 to 0) := (others => '0');
    variable r1792 : std_logic_vector(0 to 0) := (others => '0');
    variable r1791 : std_logic_vector(0 to 0) := (others => '0');
    variable r1790 : std_logic_vector(0 to 0) := (others => '0');
    variable r1789 : std_logic_vector(0 to 0) := (others => '0');
    variable r1788 : std_logic_vector(0 to 0) := (others => '0');
    variable r1787 : std_logic_vector(0 to 0) := (others => '0');
    variable r1786 : std_logic_vector(0 to 0) := (others => '0');
    variable r1785 : std_logic_vector(0 to 0) := (others => '0');
    variable r1784 : std_logic_vector(0 to 0) := (others => '0');
    variable r1783 : std_logic_vector(0 to 0) := (others => '0');
    variable r1782 : std_logic_vector(0 to 0) := (others => '0');
    variable r1781 : std_logic_vector(0 to 0) := (others => '0');
    variable r1780 : std_logic_vector(0 to 0) := (others => '0');
    variable r1779 : std_logic_vector(0 to 0) := (others => '0');
    variable r1778 : std_logic_vector(0 to 0) := (others => '0');
    variable r1777 : std_logic_vector(0 to 0) := (others => '0');
    variable r1776 : std_logic_vector(0 to 0) := (others => '0');
    variable r1775 : std_logic_vector(0 to 0) := (others => '0');
    variable r1774 : std_logic_vector(0 to 0) := (others => '0');
    variable r1773 : std_logic_vector(0 to 0) := (others => '0');
    variable r1772 : std_logic_vector(0 to 0) := (others => '0');
    variable r1771 : std_logic_vector(0 to 0) := (others => '0');
    variable r1770 : std_logic_vector(0 to 0) := (others => '0');
    variable r1769 : std_logic_vector(0 to 0) := (others => '0');
    variable r1768 : std_logic_vector(0 to 0) := (others => '0');
    variable r1767 : std_logic_vector(0 to 0) := (others => '0');
    variable r1766 : std_logic_vector(0 to 0) := (others => '0');
    variable r1765 : std_logic_vector(0 to 0) := (others => '0');
    variable r1764 : std_logic_vector(0 to 0) := (others => '0');
    variable r1763 : std_logic_vector(0 to 0) := (others => '0');
    variable r1762 : std_logic_vector(0 to 0) := (others => '0');
    variable r1761 : std_logic_vector(0 to 0) := (others => '0');
    variable r1760 : std_logic_vector(0 to 0) := (others => '0');
    variable r1759 : std_logic_vector(0 to 0) := (others => '0');
    variable r1758 : std_logic_vector(0 to 0) := (others => '0');
    variable r1757 : std_logic_vector(0 to 0) := (others => '0');
    variable r1756 : std_logic_vector(0 to 0) := (others => '0');
    variable r1755 : std_logic_vector(0 to 0) := (others => '0');
    variable r1754 : std_logic_vector(0 to 0) := (others => '0');
    variable r1753 : std_logic_vector(0 to 0) := (others => '0');
    variable r1752 : std_logic_vector(0 to 0) := (others => '0');
    variable r1751 : std_logic_vector(0 to 0) := (others => '0');
    variable r1750 : std_logic_vector(0 to 0) := (others => '0');
    variable r1749 : std_logic_vector(0 to 0) := (others => '0');
    variable r1748 : std_logic_vector(0 to 0) := (others => '0');
    variable r1747 : std_logic_vector(0 to 0) := (others => '0');
    variable r1746 : std_logic_vector(0 to 0) := (others => '0');
    variable r1745 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r1746 := "0";
    null;
    r1747 := (r1746);
    r1748 := "1";
    null;
    r1749 := (r1748);
    r1750 := "1";
    null;
    r1751 := (r1750);
    r1752 := "1";
    null;
    r1753 := (r1752);
    r1754 := "0";
    null;
    r1755 := (r1754);
    r1756 := "0";
    null;
    r1757 := (r1756);
    r1758 := "0";
    null;
    r1759 := (r1758);
    r1760 := "1";
    null;
    r1761 := (r1760);
    r1762 := "0";
    null;
    r1763 := (r1762);
    r1764 := "0";
    null;
    r1765 := (r1764);
    r1766 := "1";
    null;
    r1767 := (r1766);
    r1768 := "1";
    null;
    r1769 := (r1768);
    r1770 := "0";
    null;
    r1771 := (r1770);
    r1772 := "1";
    null;
    r1773 := (r1772);
    r1774 := "1";
    null;
    r1775 := (r1774);
    r1776 := "1";
    null;
    r1777 := (r1776);
    r1778 := "0";
    null;
    r1779 := (r1778);
    r1780 := "1";
    null;
    r1781 := (r1780);
    r1782 := "0";
    null;
    r1783 := (r1782);
    r1784 := "0";
    null;
    r1785 := (r1784);
    r1786 := "0";
    null;
    r1787 := (r1786);
    r1788 := "1";
    null;
    r1789 := (r1788);
    r1790 := "0";
    null;
    r1791 := (r1790);
    r1792 := "0";
    null;
    r1793 := (r1792);
    r1794 := "1";
    null;
    r1795 := (r1794);
    r1796 := "0";
    null;
    r1797 := (r1796);
    r1798 := "0";
    null;
    r1799 := (r1798);
    r1800 := "1";
    null;
    r1801 := (r1800);
    r1802 := "0";
    null;
    r1803 := (r1802);
    r1804 := "0";
    null;
    r1805 := (r1804);
    r1806 := "0";
    null;
    r1807 := (r1806);
    r1808 := "1";
    null;
    r1809 := (r1808);
    r1745 := (r1747 & r1749 & r1751 & r1753 & r1755 & r1757 & r1759 & r1761 & r1763 & r1765 & r1767 & r1769 & r1771 & r1773 & r1775 & r1777 & r1779 & r1781 & r1783 & r1785 & r1787 & r1789 & r1791 & r1793 & r1795 & r1797 & r1799 & r1801 & r1803 & r1805 & r1807 & r1809);
    return r1745;
  end rewire_MetaprogrammingRW.w71374491_1744;
  function rewire_MetaprogrammingRW.w428a2f98_1675 return std_logic_vector
  is
    variable r1740 : std_logic_vector(0 to 0) := (others => '0');
    variable r1739 : std_logic_vector(0 to 0) := (others => '0');
    variable r1738 : std_logic_vector(0 to 0) := (others => '0');
    variable r1737 : std_logic_vector(0 to 0) := (others => '0');
    variable r1736 : std_logic_vector(0 to 0) := (others => '0');
    variable r1735 : std_logic_vector(0 to 0) := (others => '0');
    variable r1734 : std_logic_vector(0 to 0) := (others => '0');
    variable r1733 : std_logic_vector(0 to 0) := (others => '0');
    variable r1732 : std_logic_vector(0 to 0) := (others => '0');
    variable r1731 : std_logic_vector(0 to 0) := (others => '0');
    variable r1730 : std_logic_vector(0 to 0) := (others => '0');
    variable r1729 : std_logic_vector(0 to 0) := (others => '0');
    variable r1728 : std_logic_vector(0 to 0) := (others => '0');
    variable r1727 : std_logic_vector(0 to 0) := (others => '0');
    variable r1726 : std_logic_vector(0 to 0) := (others => '0');
    variable r1725 : std_logic_vector(0 to 0) := (others => '0');
    variable r1724 : std_logic_vector(0 to 0) := (others => '0');
    variable r1723 : std_logic_vector(0 to 0) := (others => '0');
    variable r1722 : std_logic_vector(0 to 0) := (others => '0');
    variable r1721 : std_logic_vector(0 to 0) := (others => '0');
    variable r1720 : std_logic_vector(0 to 0) := (others => '0');
    variable r1719 : std_logic_vector(0 to 0) := (others => '0');
    variable r1718 : std_logic_vector(0 to 0) := (others => '0');
    variable r1717 : std_logic_vector(0 to 0) := (others => '0');
    variable r1716 : std_logic_vector(0 to 0) := (others => '0');
    variable r1715 : std_logic_vector(0 to 0) := (others => '0');
    variable r1714 : std_logic_vector(0 to 0) := (others => '0');
    variable r1713 : std_logic_vector(0 to 0) := (others => '0');
    variable r1712 : std_logic_vector(0 to 0) := (others => '0');
    variable r1711 : std_logic_vector(0 to 0) := (others => '0');
    variable r1710 : std_logic_vector(0 to 0) := (others => '0');
    variable r1709 : std_logic_vector(0 to 0) := (others => '0');
    variable r1708 : std_logic_vector(0 to 0) := (others => '0');
    variable r1707 : std_logic_vector(0 to 0) := (others => '0');
    variable r1706 : std_logic_vector(0 to 0) := (others => '0');
    variable r1705 : std_logic_vector(0 to 0) := (others => '0');
    variable r1704 : std_logic_vector(0 to 0) := (others => '0');
    variable r1703 : std_logic_vector(0 to 0) := (others => '0');
    variable r1702 : std_logic_vector(0 to 0) := (others => '0');
    variable r1701 : std_logic_vector(0 to 0) := (others => '0');
    variable r1700 : std_logic_vector(0 to 0) := (others => '0');
    variable r1699 : std_logic_vector(0 to 0) := (others => '0');
    variable r1698 : std_logic_vector(0 to 0) := (others => '0');
    variable r1697 : std_logic_vector(0 to 0) := (others => '0');
    variable r1696 : std_logic_vector(0 to 0) := (others => '0');
    variable r1695 : std_logic_vector(0 to 0) := (others => '0');
    variable r1694 : std_logic_vector(0 to 0) := (others => '0');
    variable r1693 : std_logic_vector(0 to 0) := (others => '0');
    variable r1692 : std_logic_vector(0 to 0) := (others => '0');
    variable r1691 : std_logic_vector(0 to 0) := (others => '0');
    variable r1690 : std_logic_vector(0 to 0) := (others => '0');
    variable r1689 : std_logic_vector(0 to 0) := (others => '0');
    variable r1688 : std_logic_vector(0 to 0) := (others => '0');
    variable r1687 : std_logic_vector(0 to 0) := (others => '0');
    variable r1686 : std_logic_vector(0 to 0) := (others => '0');
    variable r1685 : std_logic_vector(0 to 0) := (others => '0');
    variable r1684 : std_logic_vector(0 to 0) := (others => '0');
    variable r1683 : std_logic_vector(0 to 0) := (others => '0');
    variable r1682 : std_logic_vector(0 to 0) := (others => '0');
    variable r1681 : std_logic_vector(0 to 0) := (others => '0');
    variable r1680 : std_logic_vector(0 to 0) := (others => '0');
    variable r1679 : std_logic_vector(0 to 0) := (others => '0');
    variable r1678 : std_logic_vector(0 to 0) := (others => '0');
    variable r1677 : std_logic_vector(0 to 0) := (others => '0');
    variable r1676 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r1677 := "0";
    null;
    r1678 := (r1677);
    r1679 := "1";
    null;
    r1680 := (r1679);
    r1681 := "0";
    null;
    r1682 := (r1681);
    r1683 := "0";
    null;
    r1684 := (r1683);
    r1685 := "0";
    null;
    r1686 := (r1685);
    r1687 := "0";
    null;
    r1688 := (r1687);
    r1689 := "1";
    null;
    r1690 := (r1689);
    r1691 := "0";
    null;
    r1692 := (r1691);
    r1693 := "1";
    null;
    r1694 := (r1693);
    r1695 := "0";
    null;
    r1696 := (r1695);
    r1697 := "0";
    null;
    r1698 := (r1697);
    r1699 := "0";
    null;
    r1700 := (r1699);
    r1701 := "1";
    null;
    r1702 := (r1701);
    r1703 := "0";
    null;
    r1704 := (r1703);
    r1705 := "1";
    null;
    r1706 := (r1705);
    r1707 := "0";
    null;
    r1708 := (r1707);
    r1709 := "0";
    null;
    r1710 := (r1709);
    r1711 := "0";
    null;
    r1712 := (r1711);
    r1713 := "1";
    null;
    r1714 := (r1713);
    r1715 := "0";
    null;
    r1716 := (r1715);
    r1717 := "1";
    null;
    r1718 := (r1717);
    r1719 := "1";
    null;
    r1720 := (r1719);
    r1721 := "1";
    null;
    r1722 := (r1721);
    r1723 := "1";
    null;
    r1724 := (r1723);
    r1725 := "1";
    null;
    r1726 := (r1725);
    r1727 := "0";
    null;
    r1728 := (r1727);
    r1729 := "0";
    null;
    r1730 := (r1729);
    r1731 := "1";
    null;
    r1732 := (r1731);
    r1733 := "1";
    null;
    r1734 := (r1733);
    r1735 := "0";
    null;
    r1736 := (r1735);
    r1737 := "0";
    null;
    r1738 := (r1737);
    r1739 := "0";
    null;
    r1740 := (r1739);
    r1676 := (r1678 & r1680 & r1682 & r1684 & r1686 & r1688 & r1690 & r1692 & r1694 & r1696 & r1698 & r1700 & r1702 & r1704 & r1706 & r1708 & r1710 & r1712 & r1714 & r1716 & r1718 & r1720 & r1722 & r1724 & r1726 & r1728 & r1730 & r1732 & r1734 & r1736 & r1738 & r1740);
    return r1676;
  end rewire_MetaprogrammingRW.w428a2f98_1675;
  function rewire_Main.step256_1171(r1172 : std_logic_vector ; r1173 : std_logic_vector ; r1174 : std_logic_vector) return std_logic_vector
  is
    variable r1670 : std_logic_vector(0 to 31) := (others => '0');
    variable r1669 : std_logic_vector(0 to 31) := (others => '0');
    variable r1668 : std_logic_vector(0 to 31) := (others => '0');
    variable r1667 : std_logic_vector(0 to 31) := (others => '0');
    variable r1666 : std_logic_vector(0 to 31) := (others => '0');
    variable r1665 : std_logic_vector(0 to 31) := (others => '0');
    variable r1664 : std_logic_vector(0 to 31) := (others => '0');
    variable r1663 : std_logic_vector(0 to 31) := (others => '0');
    variable r1662 : std_logic_vector(0 to 31) := (others => '0');
    variable r1661 : std_logic_vector(0 to 31) := (others => '0');
    variable r1655 : std_logic_vector(0 to 31) := (others => '0');
    variable r1654 : std_logic_vector(0 to 31) := (others => '0');
    variable r1653 : std_logic_vector(0 to 31) := (others => '0');
    variable r1651 : std_logic_vector(0 to 31) := (others => '0');
    variable r1435 : std_logic_vector(0 to 31) := (others => '0');
    variable r1433 : std_logic_vector(0 to 31) := (others => '0');
    variable r1432 : std_logic_vector(0 to 31) := (others => '0');
    variable r1431 : std_logic_vector(0 to 31) := (others => '0');
    variable r1430 : std_logic_vector(0 to 31) := (others => '0');
    variable r1429 : std_logic_vector(0 to 31) := (others => '0');
    variable r1424 : std_logic_vector(0 to 31) := (others => '0');
    variable r1423 : std_logic_vector(0 to 31) := (others => '0');
    variable r1422 : std_logic_vector(0 to 31) := (others => '0');
    variable r1420 : std_logic_vector(0 to 31) := (others => '0');
    variable r1204 : std_logic_vector(0 to 31) := (others => '0');
    variable r1202 : std_logic_vector(0 to 255) := (others => '0');
    variable b1201 : boolean := false;
    variable b1200 : boolean := false;
    variable b1199 : boolean := false;
    variable b1198 : boolean := false;
    variable b1197 : boolean := false;
    variable b1196 : boolean := false;
    variable b1195 : boolean := false;
    variable b1194 : boolean := false;
    variable b1193 : boolean := false;
    variable b1192 : boolean := false;
    variable r1191 : std_logic_vector(0 to 31) := (others => '0');
    variable r1190 : std_logic_vector(0 to 31) := (others => '0');
    variable r1189 : std_logic_vector(0 to 31) := (others => '0');
    variable r1188 : std_logic_vector(0 to 31) := (others => '0');
    variable r1187 : std_logic_vector(0 to 31) := (others => '0');
    variable r1186 : std_logic_vector(0 to 31) := (others => '0');
    variable r1185 : std_logic_vector(0 to 31) := (others => '0');
    variable r1184 : std_logic_vector(0 to 31) := (others => '0');
    variable b1183 : boolean := false;
    variable b1182 : boolean := false;
    variable b1181 : boolean := false;
    variable r1180 : std_logic_vector(0 to 255) := (others => '0');
    variable r1179 : std_logic_vector(0 to 31) := (others => '0');
    variable r1178 : std_logic_vector(0 to 31) := (others => '0');
    variable b1177 : boolean := false;
    variable r1176 : std_logic_vector(0 to 255) := (others => '0');
    variable r1175 : std_logic_vector(0 to 319) := (others => '0');
  begin
    null;
    null;
    null;
    null;
    null;
    r1175 := (r1172 & r1173 & r1174);
    b1177 := true;
    r1178 := r1175(0 to 31);
    r1179 := r1175(32 to 63);
    r1180 := r1175(64 to 319);
    b1181 := true;
    b1182 := true;
    b1183 := true;
    r1184 := r1180(0 to 31);
    r1185 := r1180(32 to 63);
    r1186 := r1180(64 to 95);
    r1187 := r1180(96 to 127);
    r1188 := r1180(128 to 159);
    r1189 := r1180(160 to 191);
    r1190 := r1180(192 to 223);
    r1191 := r1180(224 to 255);
    b1192 := true;
    b1193 := true;
    b1194 := true;
    b1195 := true;
    b1196 := true;
    b1197 := true;
    b1198 := true;
    b1199 := true;
    b1200 := (b1183 AND (b1192 AND (b1193 AND (b1194 AND (b1195 AND (b1196 AND (b1197 AND (b1198 AND b1199))))))));
    b1201 := (b1177 AND (b1181 AND (b1182 AND b1200)));
    null;
    null;
    null;
    null;
    r1420 := rewire_Main.bigsigma1_1203(r1188);
    null;
    null;
    null;
    r1429 := rewire_Main.ch_1421(r1188,r1189,r1190);
    r1430 := w32Plus(r1420,r1429);
    null;
    null;
    r1431 := w32Plus(r1178,r1179);
    r1432 := w32Plus(r1430,r1431);
    r1433 := w32Plus(r1191,r1432);
    null;
    r1651 := rewire_Main.bigsigma0_1434(r1184);
    null;
    null;
    null;
    r1661 := rewire_Main.maj_1652(r1184,r1185,r1186);
    r1662 := w32Plus(r1651,r1661);
    r1663 := w32Plus(r1433,r1662);
    null;
    null;
    null;
    null;
    null;
    null;
    r1664 := rewire_Main.bigsigma1_1203(r1188);
    null;
    null;
    null;
    r1665 := rewire_Main.ch_1421(r1188,r1189,r1190);
    r1666 := w32Plus(r1664,r1665);
    null;
    null;
    r1667 := w32Plus(r1178,r1179);
    r1668 := w32Plus(r1666,r1667);
    r1669 := w32Plus(r1191,r1668);
    r1670 := w32Plus(r1187,r1669);
    null;
    null;
    null;
    r1202 := (r1663 & r1184 & r1185 & r1186 & r1670 & r1188 & r1189 & r1190);
    r1176 := r1202;
    return r1176;
  end rewire_Main.step256_1171;
  function rewire_Main.maj_1652(r1653 : std_logic_vector ; r1654 : std_logic_vector ; r1655 : std_logic_vector) return std_logic_vector
  is
    variable r1660 : std_logic_vector(0 to 31) := (others => '0');
    variable r1659 : std_logic_vector(0 to 31) := (others => '0');
    variable r1658 : std_logic_vector(0 to 31) := (others => '0');
    variable r1657 : std_logic_vector(0 to 31) := (others => '0');
    variable r1656 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r1656 := w32And(r1653,r1654);
    null;
    null;
    r1657 := w32And(r1653,r1655);
    r1658 := w32Xor(r1656,r1657);
    null;
    null;
    r1659 := w32And(r1654,r1655);
    r1660 := w32Xor(r1658,r1659);
    return r1660;
  end rewire_Main.maj_1652;
  function rewire_Main.bigsigma0_1434(r1435 : std_logic_vector) return std_logic_vector
  is
    variable r1650 : std_logic_vector(0 to 31) := (others => '0');
    variable r1649 : std_logic_vector(0 to 31) := (others => '0');
    variable r1580 : std_logic_vector(0 to 31) := (others => '0');
    variable r1578 : std_logic_vector(0 to 31) := (others => '0');
    variable r1577 : std_logic_vector(0 to 31) := (others => '0');
    variable r1508 : std_logic_vector(0 to 31) := (others => '0');
    variable r1506 : std_logic_vector(0 to 31) := (others => '0');
    variable r1437 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    r1506 := rewire_RWPrelude.rotateR2_1436(r1435);
    null;
    r1577 := rewire_RWPrelude.rotateR13_1507(r1435);
    r1578 := w32Xor(r1506,r1577);
    null;
    r1649 := rewire_RWPrelude.rotateR22_1579(r1435);
    r1650 := w32Xor(r1578,r1649);
    return r1650;
  end rewire_Main.bigsigma0_1434;
  function rewire_RWPrelude.rotateR22_1579(r1580 : std_logic_vector) return std_logic_vector
  is
    variable r1648 : std_logic_vector(0 to 31) := (others => '0');
    variable b1647 : boolean := false;
    variable b1646 : boolean := false;
    variable b1645 : boolean := false;
    variable b1644 : boolean := false;
    variable b1643 : boolean := false;
    variable b1642 : boolean := false;
    variable b1641 : boolean := false;
    variable b1640 : boolean := false;
    variable b1639 : boolean := false;
    variable b1638 : boolean := false;
    variable b1637 : boolean := false;
    variable b1636 : boolean := false;
    variable b1635 : boolean := false;
    variable b1634 : boolean := false;
    variable b1633 : boolean := false;
    variable b1632 : boolean := false;
    variable b1631 : boolean := false;
    variable b1630 : boolean := false;
    variable b1629 : boolean := false;
    variable b1628 : boolean := false;
    variable b1627 : boolean := false;
    variable b1626 : boolean := false;
    variable b1625 : boolean := false;
    variable b1624 : boolean := false;
    variable b1623 : boolean := false;
    variable b1622 : boolean := false;
    variable b1621 : boolean := false;
    variable b1620 : boolean := false;
    variable b1619 : boolean := false;
    variable b1618 : boolean := false;
    variable b1617 : boolean := false;
    variable b1616 : boolean := false;
    variable b1615 : boolean := false;
    variable r1614 : std_logic_vector(0 to 0) := (others => '0');
    variable r1613 : std_logic_vector(0 to 0) := (others => '0');
    variable r1612 : std_logic_vector(0 to 0) := (others => '0');
    variable r1611 : std_logic_vector(0 to 0) := (others => '0');
    variable r1610 : std_logic_vector(0 to 0) := (others => '0');
    variable r1609 : std_logic_vector(0 to 0) := (others => '0');
    variable r1608 : std_logic_vector(0 to 0) := (others => '0');
    variable r1607 : std_logic_vector(0 to 0) := (others => '0');
    variable r1606 : std_logic_vector(0 to 0) := (others => '0');
    variable r1605 : std_logic_vector(0 to 0) := (others => '0');
    variable r1604 : std_logic_vector(0 to 0) := (others => '0');
    variable r1603 : std_logic_vector(0 to 0) := (others => '0');
    variable r1602 : std_logic_vector(0 to 0) := (others => '0');
    variable r1601 : std_logic_vector(0 to 0) := (others => '0');
    variable r1600 : std_logic_vector(0 to 0) := (others => '0');
    variable r1599 : std_logic_vector(0 to 0) := (others => '0');
    variable r1598 : std_logic_vector(0 to 0) := (others => '0');
    variable r1597 : std_logic_vector(0 to 0) := (others => '0');
    variable r1596 : std_logic_vector(0 to 0) := (others => '0');
    variable r1595 : std_logic_vector(0 to 0) := (others => '0');
    variable r1594 : std_logic_vector(0 to 0) := (others => '0');
    variable r1593 : std_logic_vector(0 to 0) := (others => '0');
    variable r1592 : std_logic_vector(0 to 0) := (others => '0');
    variable r1591 : std_logic_vector(0 to 0) := (others => '0');
    variable r1590 : std_logic_vector(0 to 0) := (others => '0');
    variable r1589 : std_logic_vector(0 to 0) := (others => '0');
    variable r1588 : std_logic_vector(0 to 0) := (others => '0');
    variable r1587 : std_logic_vector(0 to 0) := (others => '0');
    variable r1586 : std_logic_vector(0 to 0) := (others => '0');
    variable r1585 : std_logic_vector(0 to 0) := (others => '0');
    variable r1584 : std_logic_vector(0 to 0) := (others => '0');
    variable r1583 : std_logic_vector(0 to 0) := (others => '0');
    variable b1582 : boolean := false;
    variable r1581 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    b1582 := true;
    r1583 := r1580(0 to 0);
    r1584 := r1580(1 to 1);
    r1585 := r1580(2 to 2);
    r1586 := r1580(3 to 3);
    r1587 := r1580(4 to 4);
    r1588 := r1580(5 to 5);
    r1589 := r1580(6 to 6);
    r1590 := r1580(7 to 7);
    r1591 := r1580(8 to 8);
    r1592 := r1580(9 to 9);
    r1593 := r1580(10 to 10);
    r1594 := r1580(11 to 11);
    r1595 := r1580(12 to 12);
    r1596 := r1580(13 to 13);
    r1597 := r1580(14 to 14);
    r1598 := r1580(15 to 15);
    r1599 := r1580(16 to 16);
    r1600 := r1580(17 to 17);
    r1601 := r1580(18 to 18);
    r1602 := r1580(19 to 19);
    r1603 := r1580(20 to 20);
    r1604 := r1580(21 to 21);
    r1605 := r1580(22 to 22);
    r1606 := r1580(23 to 23);
    r1607 := r1580(24 to 24);
    r1608 := r1580(25 to 25);
    r1609 := r1580(26 to 26);
    r1610 := r1580(27 to 27);
    r1611 := r1580(28 to 28);
    r1612 := r1580(29 to 29);
    r1613 := r1580(30 to 30);
    r1614 := r1580(31 to 31);
    b1615 := true;
    b1616 := true;
    b1617 := true;
    b1618 := true;
    b1619 := true;
    b1620 := true;
    b1621 := true;
    b1622 := true;
    b1623 := true;
    b1624 := true;
    b1625 := true;
    b1626 := true;
    b1627 := true;
    b1628 := true;
    b1629 := true;
    b1630 := true;
    b1631 := true;
    b1632 := true;
    b1633 := true;
    b1634 := true;
    b1635 := true;
    b1636 := true;
    b1637 := true;
    b1638 := true;
    b1639 := true;
    b1640 := true;
    b1641 := true;
    b1642 := true;
    b1643 := true;
    b1644 := true;
    b1645 := true;
    b1646 := true;
    b1647 := (b1582 AND (b1615 AND (b1616 AND (b1617 AND (b1618 AND (b1619 AND (b1620 AND (b1621 AND (b1622 AND (b1623 AND (b1624 AND (b1625 AND (b1626 AND (b1627 AND (b1628 AND (b1629 AND (b1630 AND (b1631 AND (b1632 AND (b1633 AND (b1634 AND (b1635 AND (b1636 AND (b1637 AND (b1638 AND (b1639 AND (b1640 AND (b1641 AND (b1642 AND (b1643 AND (b1644 AND (b1645 AND b1646))))))))))))))))))))))))))))))));
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    r1648 := (r1593 & r1594 & r1595 & r1596 & r1597 & r1598 & r1599 & r1600 & r1601 & r1602 & r1603 & r1604 & r1605 & r1606 & r1607 & r1608 & r1609 & r1610 & r1611 & r1612 & r1613 & r1614 & r1583 & r1584 & r1585 & r1586 & r1587 & r1588 & r1589 & r1590 & r1591 & r1592);
    r1581 := r1648;
    return r1581;
  end rewire_RWPrelude.rotateR22_1579;
  function rewire_RWPrelude.rotateR13_1507(r1508 : std_logic_vector) return std_logic_vector
  is
    variable r1576 : std_logic_vector(0 to 31) := (others => '0');
    variable b1575 : boolean := false;
    variable b1574 : boolean := false;
    variable b1573 : boolean := false;
    variable b1572 : boolean := false;
    variable b1571 : boolean := false;
    variable b1570 : boolean := false;
    variable b1569 : boolean := false;
    variable b1568 : boolean := false;
    variable b1567 : boolean := false;
    variable b1566 : boolean := false;
    variable b1565 : boolean := false;
    variable b1564 : boolean := false;
    variable b1563 : boolean := false;
    variable b1562 : boolean := false;
    variable b1561 : boolean := false;
    variable b1560 : boolean := false;
    variable b1559 : boolean := false;
    variable b1558 : boolean := false;
    variable b1557 : boolean := false;
    variable b1556 : boolean := false;
    variable b1555 : boolean := false;
    variable b1554 : boolean := false;
    variable b1553 : boolean := false;
    variable b1552 : boolean := false;
    variable b1551 : boolean := false;
    variable b1550 : boolean := false;
    variable b1549 : boolean := false;
    variable b1548 : boolean := false;
    variable b1547 : boolean := false;
    variable b1546 : boolean := false;
    variable b1545 : boolean := false;
    variable b1544 : boolean := false;
    variable b1543 : boolean := false;
    variable r1542 : std_logic_vector(0 to 0) := (others => '0');
    variable r1541 : std_logic_vector(0 to 0) := (others => '0');
    variable r1540 : std_logic_vector(0 to 0) := (others => '0');
    variable r1539 : std_logic_vector(0 to 0) := (others => '0');
    variable r1538 : std_logic_vector(0 to 0) := (others => '0');
    variable r1537 : std_logic_vector(0 to 0) := (others => '0');
    variable r1536 : std_logic_vector(0 to 0) := (others => '0');
    variable r1535 : std_logic_vector(0 to 0) := (others => '0');
    variable r1534 : std_logic_vector(0 to 0) := (others => '0');
    variable r1533 : std_logic_vector(0 to 0) := (others => '0');
    variable r1532 : std_logic_vector(0 to 0) := (others => '0');
    variable r1531 : std_logic_vector(0 to 0) := (others => '0');
    variable r1530 : std_logic_vector(0 to 0) := (others => '0');
    variable r1529 : std_logic_vector(0 to 0) := (others => '0');
    variable r1528 : std_logic_vector(0 to 0) := (others => '0');
    variable r1527 : std_logic_vector(0 to 0) := (others => '0');
    variable r1526 : std_logic_vector(0 to 0) := (others => '0');
    variable r1525 : std_logic_vector(0 to 0) := (others => '0');
    variable r1524 : std_logic_vector(0 to 0) := (others => '0');
    variable r1523 : std_logic_vector(0 to 0) := (others => '0');
    variable r1522 : std_logic_vector(0 to 0) := (others => '0');
    variable r1521 : std_logic_vector(0 to 0) := (others => '0');
    variable r1520 : std_logic_vector(0 to 0) := (others => '0');
    variable r1519 : std_logic_vector(0 to 0) := (others => '0');
    variable r1518 : std_logic_vector(0 to 0) := (others => '0');
    variable r1517 : std_logic_vector(0 to 0) := (others => '0');
    variable r1516 : std_logic_vector(0 to 0) := (others => '0');
    variable r1515 : std_logic_vector(0 to 0) := (others => '0');
    variable r1514 : std_logic_vector(0 to 0) := (others => '0');
    variable r1513 : std_logic_vector(0 to 0) := (others => '0');
    variable r1512 : std_logic_vector(0 to 0) := (others => '0');
    variable r1511 : std_logic_vector(0 to 0) := (others => '0');
    variable b1510 : boolean := false;
    variable r1509 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    b1510 := true;
    r1511 := r1508(0 to 0);
    r1512 := r1508(1 to 1);
    r1513 := r1508(2 to 2);
    r1514 := r1508(3 to 3);
    r1515 := r1508(4 to 4);
    r1516 := r1508(5 to 5);
    r1517 := r1508(6 to 6);
    r1518 := r1508(7 to 7);
    r1519 := r1508(8 to 8);
    r1520 := r1508(9 to 9);
    r1521 := r1508(10 to 10);
    r1522 := r1508(11 to 11);
    r1523 := r1508(12 to 12);
    r1524 := r1508(13 to 13);
    r1525 := r1508(14 to 14);
    r1526 := r1508(15 to 15);
    r1527 := r1508(16 to 16);
    r1528 := r1508(17 to 17);
    r1529 := r1508(18 to 18);
    r1530 := r1508(19 to 19);
    r1531 := r1508(20 to 20);
    r1532 := r1508(21 to 21);
    r1533 := r1508(22 to 22);
    r1534 := r1508(23 to 23);
    r1535 := r1508(24 to 24);
    r1536 := r1508(25 to 25);
    r1537 := r1508(26 to 26);
    r1538 := r1508(27 to 27);
    r1539 := r1508(28 to 28);
    r1540 := r1508(29 to 29);
    r1541 := r1508(30 to 30);
    r1542 := r1508(31 to 31);
    b1543 := true;
    b1544 := true;
    b1545 := true;
    b1546 := true;
    b1547 := true;
    b1548 := true;
    b1549 := true;
    b1550 := true;
    b1551 := true;
    b1552 := true;
    b1553 := true;
    b1554 := true;
    b1555 := true;
    b1556 := true;
    b1557 := true;
    b1558 := true;
    b1559 := true;
    b1560 := true;
    b1561 := true;
    b1562 := true;
    b1563 := true;
    b1564 := true;
    b1565 := true;
    b1566 := true;
    b1567 := true;
    b1568 := true;
    b1569 := true;
    b1570 := true;
    b1571 := true;
    b1572 := true;
    b1573 := true;
    b1574 := true;
    b1575 := (b1510 AND (b1543 AND (b1544 AND (b1545 AND (b1546 AND (b1547 AND (b1548 AND (b1549 AND (b1550 AND (b1551 AND (b1552 AND (b1553 AND (b1554 AND (b1555 AND (b1556 AND (b1557 AND (b1558 AND (b1559 AND (b1560 AND (b1561 AND (b1562 AND (b1563 AND (b1564 AND (b1565 AND (b1566 AND (b1567 AND (b1568 AND (b1569 AND (b1570 AND (b1571 AND (b1572 AND (b1573 AND b1574))))))))))))))))))))))))))))))));
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    r1576 := (r1530 & r1531 & r1532 & r1533 & r1534 & r1535 & r1536 & r1537 & r1538 & r1539 & r1540 & r1541 & r1542 & r1511 & r1512 & r1513 & r1514 & r1515 & r1516 & r1517 & r1518 & r1519 & r1520 & r1521 & r1522 & r1523 & r1524 & r1525 & r1526 & r1527 & r1528 & r1529);
    r1509 := r1576;
    return r1509;
  end rewire_RWPrelude.rotateR13_1507;
  function rewire_RWPrelude.rotateR2_1436(r1437 : std_logic_vector) return std_logic_vector
  is
    variable r1505 : std_logic_vector(0 to 31) := (others => '0');
    variable b1504 : boolean := false;
    variable b1503 : boolean := false;
    variable b1502 : boolean := false;
    variable b1501 : boolean := false;
    variable b1500 : boolean := false;
    variable b1499 : boolean := false;
    variable b1498 : boolean := false;
    variable b1497 : boolean := false;
    variable b1496 : boolean := false;
    variable b1495 : boolean := false;
    variable b1494 : boolean := false;
    variable b1493 : boolean := false;
    variable b1492 : boolean := false;
    variable b1491 : boolean := false;
    variable b1490 : boolean := false;
    variable b1489 : boolean := false;
    variable b1488 : boolean := false;
    variable b1487 : boolean := false;
    variable b1486 : boolean := false;
    variable b1485 : boolean := false;
    variable b1484 : boolean := false;
    variable b1483 : boolean := false;
    variable b1482 : boolean := false;
    variable b1481 : boolean := false;
    variable b1480 : boolean := false;
    variable b1479 : boolean := false;
    variable b1478 : boolean := false;
    variable b1477 : boolean := false;
    variable b1476 : boolean := false;
    variable b1475 : boolean := false;
    variable b1474 : boolean := false;
    variable b1473 : boolean := false;
    variable b1472 : boolean := false;
    variable r1471 : std_logic_vector(0 to 0) := (others => '0');
    variable r1470 : std_logic_vector(0 to 0) := (others => '0');
    variable r1469 : std_logic_vector(0 to 0) := (others => '0');
    variable r1468 : std_logic_vector(0 to 0) := (others => '0');
    variable r1467 : std_logic_vector(0 to 0) := (others => '0');
    variable r1466 : std_logic_vector(0 to 0) := (others => '0');
    variable r1465 : std_logic_vector(0 to 0) := (others => '0');
    variable r1464 : std_logic_vector(0 to 0) := (others => '0');
    variable r1463 : std_logic_vector(0 to 0) := (others => '0');
    variable r1462 : std_logic_vector(0 to 0) := (others => '0');
    variable r1461 : std_logic_vector(0 to 0) := (others => '0');
    variable r1460 : std_logic_vector(0 to 0) := (others => '0');
    variable r1459 : std_logic_vector(0 to 0) := (others => '0');
    variable r1458 : std_logic_vector(0 to 0) := (others => '0');
    variable r1457 : std_logic_vector(0 to 0) := (others => '0');
    variable r1456 : std_logic_vector(0 to 0) := (others => '0');
    variable r1455 : std_logic_vector(0 to 0) := (others => '0');
    variable r1454 : std_logic_vector(0 to 0) := (others => '0');
    variable r1453 : std_logic_vector(0 to 0) := (others => '0');
    variable r1452 : std_logic_vector(0 to 0) := (others => '0');
    variable r1451 : std_logic_vector(0 to 0) := (others => '0');
    variable r1450 : std_logic_vector(0 to 0) := (others => '0');
    variable r1449 : std_logic_vector(0 to 0) := (others => '0');
    variable r1448 : std_logic_vector(0 to 0) := (others => '0');
    variable r1447 : std_logic_vector(0 to 0) := (others => '0');
    variable r1446 : std_logic_vector(0 to 0) := (others => '0');
    variable r1445 : std_logic_vector(0 to 0) := (others => '0');
    variable r1444 : std_logic_vector(0 to 0) := (others => '0');
    variable r1443 : std_logic_vector(0 to 0) := (others => '0');
    variable r1442 : std_logic_vector(0 to 0) := (others => '0');
    variable r1441 : std_logic_vector(0 to 0) := (others => '0');
    variable r1440 : std_logic_vector(0 to 0) := (others => '0');
    variable b1439 : boolean := false;
    variable r1438 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    b1439 := true;
    r1440 := r1437(0 to 0);
    r1441 := r1437(1 to 1);
    r1442 := r1437(2 to 2);
    r1443 := r1437(3 to 3);
    r1444 := r1437(4 to 4);
    r1445 := r1437(5 to 5);
    r1446 := r1437(6 to 6);
    r1447 := r1437(7 to 7);
    r1448 := r1437(8 to 8);
    r1449 := r1437(9 to 9);
    r1450 := r1437(10 to 10);
    r1451 := r1437(11 to 11);
    r1452 := r1437(12 to 12);
    r1453 := r1437(13 to 13);
    r1454 := r1437(14 to 14);
    r1455 := r1437(15 to 15);
    r1456 := r1437(16 to 16);
    r1457 := r1437(17 to 17);
    r1458 := r1437(18 to 18);
    r1459 := r1437(19 to 19);
    r1460 := r1437(20 to 20);
    r1461 := r1437(21 to 21);
    r1462 := r1437(22 to 22);
    r1463 := r1437(23 to 23);
    r1464 := r1437(24 to 24);
    r1465 := r1437(25 to 25);
    r1466 := r1437(26 to 26);
    r1467 := r1437(27 to 27);
    r1468 := r1437(28 to 28);
    r1469 := r1437(29 to 29);
    r1470 := r1437(30 to 30);
    r1471 := r1437(31 to 31);
    b1472 := true;
    b1473 := true;
    b1474 := true;
    b1475 := true;
    b1476 := true;
    b1477 := true;
    b1478 := true;
    b1479 := true;
    b1480 := true;
    b1481 := true;
    b1482 := true;
    b1483 := true;
    b1484 := true;
    b1485 := true;
    b1486 := true;
    b1487 := true;
    b1488 := true;
    b1489 := true;
    b1490 := true;
    b1491 := true;
    b1492 := true;
    b1493 := true;
    b1494 := true;
    b1495 := true;
    b1496 := true;
    b1497 := true;
    b1498 := true;
    b1499 := true;
    b1500 := true;
    b1501 := true;
    b1502 := true;
    b1503 := true;
    b1504 := (b1439 AND (b1472 AND (b1473 AND (b1474 AND (b1475 AND (b1476 AND (b1477 AND (b1478 AND (b1479 AND (b1480 AND (b1481 AND (b1482 AND (b1483 AND (b1484 AND (b1485 AND (b1486 AND (b1487 AND (b1488 AND (b1489 AND (b1490 AND (b1491 AND (b1492 AND (b1493 AND (b1494 AND (b1495 AND (b1496 AND (b1497 AND (b1498 AND (b1499 AND (b1500 AND (b1501 AND (b1502 AND b1503))))))))))))))))))))))))))))))));
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    r1505 := (r1470 & r1471 & r1440 & r1441 & r1442 & r1443 & r1444 & r1445 & r1446 & r1447 & r1448 & r1449 & r1450 & r1451 & r1452 & r1453 & r1454 & r1455 & r1456 & r1457 & r1458 & r1459 & r1460 & r1461 & r1462 & r1463 & r1464 & r1465 & r1466 & r1467 & r1468 & r1469);
    r1438 := r1505;
    return r1438;
  end rewire_RWPrelude.rotateR2_1436;
  function rewire_Main.ch_1421(r1422 : std_logic_vector ; r1423 : std_logic_vector ; r1424 : std_logic_vector) return std_logic_vector
  is
    variable r1428 : std_logic_vector(0 to 31) := (others => '0');
    variable r1427 : std_logic_vector(0 to 31) := (others => '0');
    variable r1426 : std_logic_vector(0 to 31) := (others => '0');
    variable r1425 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r1425 := w32And(r1422,r1423);
    null;
    r1426 := w32Not(r1422);
    null;
    r1427 := w32And(r1426,r1424);
    r1428 := w32Xor(r1425,r1427);
    return r1428;
  end rewire_Main.ch_1421;
  function rewire_Main.bigsigma1_1203(r1204 : std_logic_vector) return std_logic_vector
  is
    variable r1419 : std_logic_vector(0 to 31) := (others => '0');
    variable r1418 : std_logic_vector(0 to 31) := (others => '0');
    variable r1349 : std_logic_vector(0 to 31) := (others => '0');
    variable r1347 : std_logic_vector(0 to 31) := (others => '0');
    variable r1346 : std_logic_vector(0 to 31) := (others => '0');
    variable r1277 : std_logic_vector(0 to 31) := (others => '0');
    variable r1275 : std_logic_vector(0 to 31) := (others => '0');
    variable r1206 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    r1275 := rewire_RWPrelude.rotateR6_1205(r1204);
    null;
    r1346 := rewire_RWPrelude.rotateR11_1276(r1204);
    r1347 := w32Xor(r1275,r1346);
    null;
    r1418 := rewire_RWPrelude.rotateR25_1348(r1204);
    r1419 := w32Xor(r1347,r1418);
    return r1419;
  end rewire_Main.bigsigma1_1203;
  function rewire_RWPrelude.rotateR25_1348(r1349 : std_logic_vector) return std_logic_vector
  is
    variable r1417 : std_logic_vector(0 to 31) := (others => '0');
    variable b1416 : boolean := false;
    variable b1415 : boolean := false;
    variable b1414 : boolean := false;
    variable b1413 : boolean := false;
    variable b1412 : boolean := false;
    variable b1411 : boolean := false;
    variable b1410 : boolean := false;
    variable b1409 : boolean := false;
    variable b1408 : boolean := false;
    variable b1407 : boolean := false;
    variable b1406 : boolean := false;
    variable b1405 : boolean := false;
    variable b1404 : boolean := false;
    variable b1403 : boolean := false;
    variable b1402 : boolean := false;
    variable b1401 : boolean := false;
    variable b1400 : boolean := false;
    variable b1399 : boolean := false;
    variable b1398 : boolean := false;
    variable b1397 : boolean := false;
    variable b1396 : boolean := false;
    variable b1395 : boolean := false;
    variable b1394 : boolean := false;
    variable b1393 : boolean := false;
    variable b1392 : boolean := false;
    variable b1391 : boolean := false;
    variable b1390 : boolean := false;
    variable b1389 : boolean := false;
    variable b1388 : boolean := false;
    variable b1387 : boolean := false;
    variable b1386 : boolean := false;
    variable b1385 : boolean := false;
    variable b1384 : boolean := false;
    variable r1383 : std_logic_vector(0 to 0) := (others => '0');
    variable r1382 : std_logic_vector(0 to 0) := (others => '0');
    variable r1381 : std_logic_vector(0 to 0) := (others => '0');
    variable r1380 : std_logic_vector(0 to 0) := (others => '0');
    variable r1379 : std_logic_vector(0 to 0) := (others => '0');
    variable r1378 : std_logic_vector(0 to 0) := (others => '0');
    variable r1377 : std_logic_vector(0 to 0) := (others => '0');
    variable r1376 : std_logic_vector(0 to 0) := (others => '0');
    variable r1375 : std_logic_vector(0 to 0) := (others => '0');
    variable r1374 : std_logic_vector(0 to 0) := (others => '0');
    variable r1373 : std_logic_vector(0 to 0) := (others => '0');
    variable r1372 : std_logic_vector(0 to 0) := (others => '0');
    variable r1371 : std_logic_vector(0 to 0) := (others => '0');
    variable r1370 : std_logic_vector(0 to 0) := (others => '0');
    variable r1369 : std_logic_vector(0 to 0) := (others => '0');
    variable r1368 : std_logic_vector(0 to 0) := (others => '0');
    variable r1367 : std_logic_vector(0 to 0) := (others => '0');
    variable r1366 : std_logic_vector(0 to 0) := (others => '0');
    variable r1365 : std_logic_vector(0 to 0) := (others => '0');
    variable r1364 : std_logic_vector(0 to 0) := (others => '0');
    variable r1363 : std_logic_vector(0 to 0) := (others => '0');
    variable r1362 : std_logic_vector(0 to 0) := (others => '0');
    variable r1361 : std_logic_vector(0 to 0) := (others => '0');
    variable r1360 : std_logic_vector(0 to 0) := (others => '0');
    variable r1359 : std_logic_vector(0 to 0) := (others => '0');
    variable r1358 : std_logic_vector(0 to 0) := (others => '0');
    variable r1357 : std_logic_vector(0 to 0) := (others => '0');
    variable r1356 : std_logic_vector(0 to 0) := (others => '0');
    variable r1355 : std_logic_vector(0 to 0) := (others => '0');
    variable r1354 : std_logic_vector(0 to 0) := (others => '0');
    variable r1353 : std_logic_vector(0 to 0) := (others => '0');
    variable r1352 : std_logic_vector(0 to 0) := (others => '0');
    variable b1351 : boolean := false;
    variable r1350 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    b1351 := true;
    r1352 := r1349(0 to 0);
    r1353 := r1349(1 to 1);
    r1354 := r1349(2 to 2);
    r1355 := r1349(3 to 3);
    r1356 := r1349(4 to 4);
    r1357 := r1349(5 to 5);
    r1358 := r1349(6 to 6);
    r1359 := r1349(7 to 7);
    r1360 := r1349(8 to 8);
    r1361 := r1349(9 to 9);
    r1362 := r1349(10 to 10);
    r1363 := r1349(11 to 11);
    r1364 := r1349(12 to 12);
    r1365 := r1349(13 to 13);
    r1366 := r1349(14 to 14);
    r1367 := r1349(15 to 15);
    r1368 := r1349(16 to 16);
    r1369 := r1349(17 to 17);
    r1370 := r1349(18 to 18);
    r1371 := r1349(19 to 19);
    r1372 := r1349(20 to 20);
    r1373 := r1349(21 to 21);
    r1374 := r1349(22 to 22);
    r1375 := r1349(23 to 23);
    r1376 := r1349(24 to 24);
    r1377 := r1349(25 to 25);
    r1378 := r1349(26 to 26);
    r1379 := r1349(27 to 27);
    r1380 := r1349(28 to 28);
    r1381 := r1349(29 to 29);
    r1382 := r1349(30 to 30);
    r1383 := r1349(31 to 31);
    b1384 := true;
    b1385 := true;
    b1386 := true;
    b1387 := true;
    b1388 := true;
    b1389 := true;
    b1390 := true;
    b1391 := true;
    b1392 := true;
    b1393 := true;
    b1394 := true;
    b1395 := true;
    b1396 := true;
    b1397 := true;
    b1398 := true;
    b1399 := true;
    b1400 := true;
    b1401 := true;
    b1402 := true;
    b1403 := true;
    b1404 := true;
    b1405 := true;
    b1406 := true;
    b1407 := true;
    b1408 := true;
    b1409 := true;
    b1410 := true;
    b1411 := true;
    b1412 := true;
    b1413 := true;
    b1414 := true;
    b1415 := true;
    b1416 := (b1351 AND (b1384 AND (b1385 AND (b1386 AND (b1387 AND (b1388 AND (b1389 AND (b1390 AND (b1391 AND (b1392 AND (b1393 AND (b1394 AND (b1395 AND (b1396 AND (b1397 AND (b1398 AND (b1399 AND (b1400 AND (b1401 AND (b1402 AND (b1403 AND (b1404 AND (b1405 AND (b1406 AND (b1407 AND (b1408 AND (b1409 AND (b1410 AND (b1411 AND (b1412 AND (b1413 AND (b1414 AND b1415))))))))))))))))))))))))))))))));
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    r1417 := (r1359 & r1360 & r1361 & r1362 & r1363 & r1364 & r1365 & r1366 & r1367 & r1368 & r1369 & r1370 & r1371 & r1372 & r1373 & r1374 & r1375 & r1376 & r1377 & r1378 & r1379 & r1380 & r1381 & r1382 & r1383 & r1352 & r1353 & r1354 & r1355 & r1356 & r1357 & r1358);
    r1350 := r1417;
    return r1350;
  end rewire_RWPrelude.rotateR25_1348;
  function rewire_RWPrelude.rotateR11_1276(r1277 : std_logic_vector) return std_logic_vector
  is
    variable r1345 : std_logic_vector(0 to 31) := (others => '0');
    variable b1344 : boolean := false;
    variable b1343 : boolean := false;
    variable b1342 : boolean := false;
    variable b1341 : boolean := false;
    variable b1340 : boolean := false;
    variable b1339 : boolean := false;
    variable b1338 : boolean := false;
    variable b1337 : boolean := false;
    variable b1336 : boolean := false;
    variable b1335 : boolean := false;
    variable b1334 : boolean := false;
    variable b1333 : boolean := false;
    variable b1332 : boolean := false;
    variable b1331 : boolean := false;
    variable b1330 : boolean := false;
    variable b1329 : boolean := false;
    variable b1328 : boolean := false;
    variable b1327 : boolean := false;
    variable b1326 : boolean := false;
    variable b1325 : boolean := false;
    variable b1324 : boolean := false;
    variable b1323 : boolean := false;
    variable b1322 : boolean := false;
    variable b1321 : boolean := false;
    variable b1320 : boolean := false;
    variable b1319 : boolean := false;
    variable b1318 : boolean := false;
    variable b1317 : boolean := false;
    variable b1316 : boolean := false;
    variable b1315 : boolean := false;
    variable b1314 : boolean := false;
    variable b1313 : boolean := false;
    variable b1312 : boolean := false;
    variable r1311 : std_logic_vector(0 to 0) := (others => '0');
    variable r1310 : std_logic_vector(0 to 0) := (others => '0');
    variable r1309 : std_logic_vector(0 to 0) := (others => '0');
    variable r1308 : std_logic_vector(0 to 0) := (others => '0');
    variable r1307 : std_logic_vector(0 to 0) := (others => '0');
    variable r1306 : std_logic_vector(0 to 0) := (others => '0');
    variable r1305 : std_logic_vector(0 to 0) := (others => '0');
    variable r1304 : std_logic_vector(0 to 0) := (others => '0');
    variable r1303 : std_logic_vector(0 to 0) := (others => '0');
    variable r1302 : std_logic_vector(0 to 0) := (others => '0');
    variable r1301 : std_logic_vector(0 to 0) := (others => '0');
    variable r1300 : std_logic_vector(0 to 0) := (others => '0');
    variable r1299 : std_logic_vector(0 to 0) := (others => '0');
    variable r1298 : std_logic_vector(0 to 0) := (others => '0');
    variable r1297 : std_logic_vector(0 to 0) := (others => '0');
    variable r1296 : std_logic_vector(0 to 0) := (others => '0');
    variable r1295 : std_logic_vector(0 to 0) := (others => '0');
    variable r1294 : std_logic_vector(0 to 0) := (others => '0');
    variable r1293 : std_logic_vector(0 to 0) := (others => '0');
    variable r1292 : std_logic_vector(0 to 0) := (others => '0');
    variable r1291 : std_logic_vector(0 to 0) := (others => '0');
    variable r1290 : std_logic_vector(0 to 0) := (others => '0');
    variable r1289 : std_logic_vector(0 to 0) := (others => '0');
    variable r1288 : std_logic_vector(0 to 0) := (others => '0');
    variable r1287 : std_logic_vector(0 to 0) := (others => '0');
    variable r1286 : std_logic_vector(0 to 0) := (others => '0');
    variable r1285 : std_logic_vector(0 to 0) := (others => '0');
    variable r1284 : std_logic_vector(0 to 0) := (others => '0');
    variable r1283 : std_logic_vector(0 to 0) := (others => '0');
    variable r1282 : std_logic_vector(0 to 0) := (others => '0');
    variable r1281 : std_logic_vector(0 to 0) := (others => '0');
    variable r1280 : std_logic_vector(0 to 0) := (others => '0');
    variable b1279 : boolean := false;
    variable r1278 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    b1279 := true;
    r1280 := r1277(0 to 0);
    r1281 := r1277(1 to 1);
    r1282 := r1277(2 to 2);
    r1283 := r1277(3 to 3);
    r1284 := r1277(4 to 4);
    r1285 := r1277(5 to 5);
    r1286 := r1277(6 to 6);
    r1287 := r1277(7 to 7);
    r1288 := r1277(8 to 8);
    r1289 := r1277(9 to 9);
    r1290 := r1277(10 to 10);
    r1291 := r1277(11 to 11);
    r1292 := r1277(12 to 12);
    r1293 := r1277(13 to 13);
    r1294 := r1277(14 to 14);
    r1295 := r1277(15 to 15);
    r1296 := r1277(16 to 16);
    r1297 := r1277(17 to 17);
    r1298 := r1277(18 to 18);
    r1299 := r1277(19 to 19);
    r1300 := r1277(20 to 20);
    r1301 := r1277(21 to 21);
    r1302 := r1277(22 to 22);
    r1303 := r1277(23 to 23);
    r1304 := r1277(24 to 24);
    r1305 := r1277(25 to 25);
    r1306 := r1277(26 to 26);
    r1307 := r1277(27 to 27);
    r1308 := r1277(28 to 28);
    r1309 := r1277(29 to 29);
    r1310 := r1277(30 to 30);
    r1311 := r1277(31 to 31);
    b1312 := true;
    b1313 := true;
    b1314 := true;
    b1315 := true;
    b1316 := true;
    b1317 := true;
    b1318 := true;
    b1319 := true;
    b1320 := true;
    b1321 := true;
    b1322 := true;
    b1323 := true;
    b1324 := true;
    b1325 := true;
    b1326 := true;
    b1327 := true;
    b1328 := true;
    b1329 := true;
    b1330 := true;
    b1331 := true;
    b1332 := true;
    b1333 := true;
    b1334 := true;
    b1335 := true;
    b1336 := true;
    b1337 := true;
    b1338 := true;
    b1339 := true;
    b1340 := true;
    b1341 := true;
    b1342 := true;
    b1343 := true;
    b1344 := (b1279 AND (b1312 AND (b1313 AND (b1314 AND (b1315 AND (b1316 AND (b1317 AND (b1318 AND (b1319 AND (b1320 AND (b1321 AND (b1322 AND (b1323 AND (b1324 AND (b1325 AND (b1326 AND (b1327 AND (b1328 AND (b1329 AND (b1330 AND (b1331 AND (b1332 AND (b1333 AND (b1334 AND (b1335 AND (b1336 AND (b1337 AND (b1338 AND (b1339 AND (b1340 AND (b1341 AND (b1342 AND b1343))))))))))))))))))))))))))))))));
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    r1345 := (r1301 & r1302 & r1303 & r1304 & r1305 & r1306 & r1307 & r1308 & r1309 & r1310 & r1311 & r1280 & r1281 & r1282 & r1283 & r1284 & r1285 & r1286 & r1287 & r1288 & r1289 & r1290 & r1291 & r1292 & r1293 & r1294 & r1295 & r1296 & r1297 & r1298 & r1299 & r1300);
    r1278 := r1345;
    return r1278;
  end rewire_RWPrelude.rotateR11_1276;
  function rewire_RWPrelude.rotateR6_1205(r1206 : std_logic_vector) return std_logic_vector
  is
    variable r1274 : std_logic_vector(0 to 31) := (others => '0');
    variable b1273 : boolean := false;
    variable b1272 : boolean := false;
    variable b1271 : boolean := false;
    variable b1270 : boolean := false;
    variable b1269 : boolean := false;
    variable b1268 : boolean := false;
    variable b1267 : boolean := false;
    variable b1266 : boolean := false;
    variable b1265 : boolean := false;
    variable b1264 : boolean := false;
    variable b1263 : boolean := false;
    variable b1262 : boolean := false;
    variable b1261 : boolean := false;
    variable b1260 : boolean := false;
    variable b1259 : boolean := false;
    variable b1258 : boolean := false;
    variable b1257 : boolean := false;
    variable b1256 : boolean := false;
    variable b1255 : boolean := false;
    variable b1254 : boolean := false;
    variable b1253 : boolean := false;
    variable b1252 : boolean := false;
    variable b1251 : boolean := false;
    variable b1250 : boolean := false;
    variable b1249 : boolean := false;
    variable b1248 : boolean := false;
    variable b1247 : boolean := false;
    variable b1246 : boolean := false;
    variable b1245 : boolean := false;
    variable b1244 : boolean := false;
    variable b1243 : boolean := false;
    variable b1242 : boolean := false;
    variable b1241 : boolean := false;
    variable r1240 : std_logic_vector(0 to 0) := (others => '0');
    variable r1239 : std_logic_vector(0 to 0) := (others => '0');
    variable r1238 : std_logic_vector(0 to 0) := (others => '0');
    variable r1237 : std_logic_vector(0 to 0) := (others => '0');
    variable r1236 : std_logic_vector(0 to 0) := (others => '0');
    variable r1235 : std_logic_vector(0 to 0) := (others => '0');
    variable r1234 : std_logic_vector(0 to 0) := (others => '0');
    variable r1233 : std_logic_vector(0 to 0) := (others => '0');
    variable r1232 : std_logic_vector(0 to 0) := (others => '0');
    variable r1231 : std_logic_vector(0 to 0) := (others => '0');
    variable r1230 : std_logic_vector(0 to 0) := (others => '0');
    variable r1229 : std_logic_vector(0 to 0) := (others => '0');
    variable r1228 : std_logic_vector(0 to 0) := (others => '0');
    variable r1227 : std_logic_vector(0 to 0) := (others => '0');
    variable r1226 : std_logic_vector(0 to 0) := (others => '0');
    variable r1225 : std_logic_vector(0 to 0) := (others => '0');
    variable r1224 : std_logic_vector(0 to 0) := (others => '0');
    variable r1223 : std_logic_vector(0 to 0) := (others => '0');
    variable r1222 : std_logic_vector(0 to 0) := (others => '0');
    variable r1221 : std_logic_vector(0 to 0) := (others => '0');
    variable r1220 : std_logic_vector(0 to 0) := (others => '0');
    variable r1219 : std_logic_vector(0 to 0) := (others => '0');
    variable r1218 : std_logic_vector(0 to 0) := (others => '0');
    variable r1217 : std_logic_vector(0 to 0) := (others => '0');
    variable r1216 : std_logic_vector(0 to 0) := (others => '0');
    variable r1215 : std_logic_vector(0 to 0) := (others => '0');
    variable r1214 : std_logic_vector(0 to 0) := (others => '0');
    variable r1213 : std_logic_vector(0 to 0) := (others => '0');
    variable r1212 : std_logic_vector(0 to 0) := (others => '0');
    variable r1211 : std_logic_vector(0 to 0) := (others => '0');
    variable r1210 : std_logic_vector(0 to 0) := (others => '0');
    variable r1209 : std_logic_vector(0 to 0) := (others => '0');
    variable b1208 : boolean := false;
    variable r1207 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    b1208 := true;
    r1209 := r1206(0 to 0);
    r1210 := r1206(1 to 1);
    r1211 := r1206(2 to 2);
    r1212 := r1206(3 to 3);
    r1213 := r1206(4 to 4);
    r1214 := r1206(5 to 5);
    r1215 := r1206(6 to 6);
    r1216 := r1206(7 to 7);
    r1217 := r1206(8 to 8);
    r1218 := r1206(9 to 9);
    r1219 := r1206(10 to 10);
    r1220 := r1206(11 to 11);
    r1221 := r1206(12 to 12);
    r1222 := r1206(13 to 13);
    r1223 := r1206(14 to 14);
    r1224 := r1206(15 to 15);
    r1225 := r1206(16 to 16);
    r1226 := r1206(17 to 17);
    r1227 := r1206(18 to 18);
    r1228 := r1206(19 to 19);
    r1229 := r1206(20 to 20);
    r1230 := r1206(21 to 21);
    r1231 := r1206(22 to 22);
    r1232 := r1206(23 to 23);
    r1233 := r1206(24 to 24);
    r1234 := r1206(25 to 25);
    r1235 := r1206(26 to 26);
    r1236 := r1206(27 to 27);
    r1237 := r1206(28 to 28);
    r1238 := r1206(29 to 29);
    r1239 := r1206(30 to 30);
    r1240 := r1206(31 to 31);
    b1241 := true;
    b1242 := true;
    b1243 := true;
    b1244 := true;
    b1245 := true;
    b1246 := true;
    b1247 := true;
    b1248 := true;
    b1249 := true;
    b1250 := true;
    b1251 := true;
    b1252 := true;
    b1253 := true;
    b1254 := true;
    b1255 := true;
    b1256 := true;
    b1257 := true;
    b1258 := true;
    b1259 := true;
    b1260 := true;
    b1261 := true;
    b1262 := true;
    b1263 := true;
    b1264 := true;
    b1265 := true;
    b1266 := true;
    b1267 := true;
    b1268 := true;
    b1269 := true;
    b1270 := true;
    b1271 := true;
    b1272 := true;
    b1273 := (b1208 AND (b1241 AND (b1242 AND (b1243 AND (b1244 AND (b1245 AND (b1246 AND (b1247 AND (b1248 AND (b1249 AND (b1250 AND (b1251 AND (b1252 AND (b1253 AND (b1254 AND (b1255 AND (b1256 AND (b1257 AND (b1258 AND (b1259 AND (b1260 AND (b1261 AND (b1262 AND (b1263 AND (b1264 AND (b1265 AND (b1266 AND (b1267 AND (b1268 AND (b1269 AND (b1270 AND (b1271 AND b1272))))))))))))))))))))))))))))))));
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    r1274 := (r1235 & r1236 & r1237 & r1238 & r1239 & r1240 & r1209 & r1210 & r1211 & r1212 & r1213 & r1214 & r1215 & r1216 & r1217 & r1218 & r1219 & r1220 & r1221 & r1222 & r1223 & r1224 & r1225 & r1226 & r1227 & r1228 & r1229 & r1230 & r1231 & r1232 & r1233 & r1234);
    r1207 := r1274;
    return r1207;
  end rewire_RWPrelude.rotateR6_1205;
  function rewire_Main.updateSched_659(r660 : std_logic_vector) return std_logic_vector
  is
    variable r1161 : std_logic_vector(0 to 31) := (others => '0');
    variable r1160 : std_logic_vector(0 to 31) := (others => '0');
    variable r1159 : std_logic_vector(0 to 31) := (others => '0');
    variable r937 : std_logic_vector(0 to 31) := (others => '0');
    variable r935 : std_logic_vector(0 to 31) := (others => '0');
    variable r934 : std_logic_vector(0 to 31) := (others => '0');
    variable r698 : std_logic_vector(0 to 31) := (others => '0');
    variable r696 : std_logic_vector(0 to 511) := (others => '0');
    variable b695 : boolean := false;
    variable b694 : boolean := false;
    variable b693 : boolean := false;
    variable b692 : boolean := false;
    variable b691 : boolean := false;
    variable b690 : boolean := false;
    variable b689 : boolean := false;
    variable b688 : boolean := false;
    variable b687 : boolean := false;
    variable b686 : boolean := false;
    variable b685 : boolean := false;
    variable b684 : boolean := false;
    variable b683 : boolean := false;
    variable b682 : boolean := false;
    variable b681 : boolean := false;
    variable b680 : boolean := false;
    variable b679 : boolean := false;
    variable r678 : std_logic_vector(0 to 31) := (others => '0');
    variable r677 : std_logic_vector(0 to 31) := (others => '0');
    variable r676 : std_logic_vector(0 to 31) := (others => '0');
    variable r675 : std_logic_vector(0 to 31) := (others => '0');
    variable r674 : std_logic_vector(0 to 31) := (others => '0');
    variable r673 : std_logic_vector(0 to 31) := (others => '0');
    variable r672 : std_logic_vector(0 to 31) := (others => '0');
    variable r671 : std_logic_vector(0 to 31) := (others => '0');
    variable r670 : std_logic_vector(0 to 31) := (others => '0');
    variable r669 : std_logic_vector(0 to 31) := (others => '0');
    variable r668 : std_logic_vector(0 to 31) := (others => '0');
    variable r667 : std_logic_vector(0 to 31) := (others => '0');
    variable r666 : std_logic_vector(0 to 31) := (others => '0');
    variable r665 : std_logic_vector(0 to 31) := (others => '0');
    variable r664 : std_logic_vector(0 to 31) := (others => '0');
    variable r663 : std_logic_vector(0 to 31) := (others => '0');
    variable b662 : boolean := false;
    variable r661 : std_logic_vector(0 to 511) := (others => '0');
  begin
    null;
    b662 := true;
    r663 := r660(0 to 31);
    r664 := r660(32 to 63);
    r665 := r660(64 to 95);
    r666 := r660(96 to 127);
    r667 := r660(128 to 159);
    r668 := r660(160 to 191);
    r669 := r660(192 to 223);
    r670 := r660(224 to 255);
    r671 := r660(256 to 287);
    r672 := r660(288 to 319);
    r673 := r660(320 to 351);
    r674 := r660(352 to 383);
    r675 := r660(384 to 415);
    r676 := r660(416 to 447);
    r677 := r660(448 to 479);
    r678 := r660(480 to 511);
    b679 := true;
    b680 := true;
    b681 := true;
    b682 := true;
    b683 := true;
    b684 := true;
    b685 := true;
    b686 := true;
    b687 := true;
    b688 := true;
    b689 := true;
    b690 := true;
    b691 := true;
    b692 := true;
    b693 := true;
    b694 := true;
    b695 := (b662 AND (b679 AND (b680 AND (b681 AND (b682 AND (b683 AND (b684 AND (b685 AND (b686 AND (b687 AND (b688 AND (b689 AND (b690 AND (b691 AND (b692 AND (b693 AND b694))))))))))))))));
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    r934 := rewire_Main.sigma1_697(r677);
    null;
    r935 := w32Plus(r934,r672);
    null;
    r1159 := rewire_Main.sigma0_936(r664);
    null;
    r1160 := w32Plus(r1159,r663);
    r1161 := w32Plus(r935,r1160);
    r696 := (r664 & r665 & r666 & r667 & r668 & r669 & r670 & r671 & r672 & r673 & r674 & r675 & r676 & r677 & r678 & r1161);
    r661 := r696;
    return r661;
  end rewire_Main.updateSched_659;
  function rewire_Main.sigma0_936(r937 : std_logic_vector) return std_logic_vector
  is
    variable r1158 : std_logic_vector(0 to 31) := (others => '0');
    variable r1157 : std_logic_vector(0 to 31) := (others => '0');
    variable r1082 : std_logic_vector(0 to 31) := (others => '0');
    variable r1080 : std_logic_vector(0 to 31) := (others => '0');
    variable r1079 : std_logic_vector(0 to 31) := (others => '0');
    variable r1010 : std_logic_vector(0 to 31) := (others => '0');
    variable r1008 : std_logic_vector(0 to 31) := (others => '0');
    variable r939 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    r1008 := rewire_RWPrelude.rotateR7_938(r937);
    null;
    r1079 := rewire_RWPrelude.rotateR18_1009(r937);
    r1080 := w32Xor(r1008,r1079);
    null;
    r1157 := rewire_RWPrelude.shiftR3_1081(r937);
    r1158 := w32Xor(r1080,r1157);
    return r1158;
  end rewire_Main.sigma0_936;
  function rewire_RWPrelude.shiftR3_1081(r1082 : std_logic_vector) return std_logic_vector
  is
    variable r1156 : std_logic_vector(0 to 0) := (others => '0');
    variable r1155 : std_logic_vector(0 to 0) := (others => '0');
    variable r1154 : std_logic_vector(0 to 0) := (others => '0');
    variable r1153 : std_logic_vector(0 to 0) := (others => '0');
    variable r1152 : std_logic_vector(0 to 0) := (others => '0');
    variable r1151 : std_logic_vector(0 to 0) := (others => '0');
    variable r1150 : std_logic_vector(0 to 31) := (others => '0');
    variable b1149 : boolean := false;
    variable b1148 : boolean := false;
    variable b1147 : boolean := false;
    variable b1146 : boolean := false;
    variable b1145 : boolean := false;
    variable b1144 : boolean := false;
    variable b1143 : boolean := false;
    variable b1142 : boolean := false;
    variable b1141 : boolean := false;
    variable b1140 : boolean := false;
    variable b1139 : boolean := false;
    variable b1138 : boolean := false;
    variable b1137 : boolean := false;
    variable b1136 : boolean := false;
    variable b1135 : boolean := false;
    variable b1134 : boolean := false;
    variable b1133 : boolean := false;
    variable b1132 : boolean := false;
    variable b1131 : boolean := false;
    variable b1130 : boolean := false;
    variable b1129 : boolean := false;
    variable b1128 : boolean := false;
    variable b1127 : boolean := false;
    variable b1126 : boolean := false;
    variable b1125 : boolean := false;
    variable b1124 : boolean := false;
    variable b1123 : boolean := false;
    variable b1122 : boolean := false;
    variable b1121 : boolean := false;
    variable b1120 : boolean := false;
    variable b1119 : boolean := false;
    variable b1118 : boolean := false;
    variable b1117 : boolean := false;
    variable r1116 : std_logic_vector(0 to 0) := (others => '0');
    variable r1115 : std_logic_vector(0 to 0) := (others => '0');
    variable r1114 : std_logic_vector(0 to 0) := (others => '0');
    variable r1113 : std_logic_vector(0 to 0) := (others => '0');
    variable r1112 : std_logic_vector(0 to 0) := (others => '0');
    variable r1111 : std_logic_vector(0 to 0) := (others => '0');
    variable r1110 : std_logic_vector(0 to 0) := (others => '0');
    variable r1109 : std_logic_vector(0 to 0) := (others => '0');
    variable r1108 : std_logic_vector(0 to 0) := (others => '0');
    variable r1107 : std_logic_vector(0 to 0) := (others => '0');
    variable r1106 : std_logic_vector(0 to 0) := (others => '0');
    variable r1105 : std_logic_vector(0 to 0) := (others => '0');
    variable r1104 : std_logic_vector(0 to 0) := (others => '0');
    variable r1103 : std_logic_vector(0 to 0) := (others => '0');
    variable r1102 : std_logic_vector(0 to 0) := (others => '0');
    variable r1101 : std_logic_vector(0 to 0) := (others => '0');
    variable r1100 : std_logic_vector(0 to 0) := (others => '0');
    variable r1099 : std_logic_vector(0 to 0) := (others => '0');
    variable r1098 : std_logic_vector(0 to 0) := (others => '0');
    variable r1097 : std_logic_vector(0 to 0) := (others => '0');
    variable r1096 : std_logic_vector(0 to 0) := (others => '0');
    variable r1095 : std_logic_vector(0 to 0) := (others => '0');
    variable r1094 : std_logic_vector(0 to 0) := (others => '0');
    variable r1093 : std_logic_vector(0 to 0) := (others => '0');
    variable r1092 : std_logic_vector(0 to 0) := (others => '0');
    variable r1091 : std_logic_vector(0 to 0) := (others => '0');
    variable r1090 : std_logic_vector(0 to 0) := (others => '0');
    variable r1089 : std_logic_vector(0 to 0) := (others => '0');
    variable r1088 : std_logic_vector(0 to 0) := (others => '0');
    variable r1087 : std_logic_vector(0 to 0) := (others => '0');
    variable r1086 : std_logic_vector(0 to 0) := (others => '0');
    variable r1085 : std_logic_vector(0 to 0) := (others => '0');
    variable b1084 : boolean := false;
    variable r1083 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    b1084 := true;
    r1085 := r1082(0 to 0);
    r1086 := r1082(1 to 1);
    r1087 := r1082(2 to 2);
    r1088 := r1082(3 to 3);
    r1089 := r1082(4 to 4);
    r1090 := r1082(5 to 5);
    r1091 := r1082(6 to 6);
    r1092 := r1082(7 to 7);
    r1093 := r1082(8 to 8);
    r1094 := r1082(9 to 9);
    r1095 := r1082(10 to 10);
    r1096 := r1082(11 to 11);
    r1097 := r1082(12 to 12);
    r1098 := r1082(13 to 13);
    r1099 := r1082(14 to 14);
    r1100 := r1082(15 to 15);
    r1101 := r1082(16 to 16);
    r1102 := r1082(17 to 17);
    r1103 := r1082(18 to 18);
    r1104 := r1082(19 to 19);
    r1105 := r1082(20 to 20);
    r1106 := r1082(21 to 21);
    r1107 := r1082(22 to 22);
    r1108 := r1082(23 to 23);
    r1109 := r1082(24 to 24);
    r1110 := r1082(25 to 25);
    r1111 := r1082(26 to 26);
    r1112 := r1082(27 to 27);
    r1113 := r1082(28 to 28);
    r1114 := r1082(29 to 29);
    r1115 := r1082(30 to 30);
    r1116 := r1082(31 to 31);
    b1117 := true;
    b1118 := true;
    b1119 := true;
    b1120 := true;
    b1121 := true;
    b1122 := true;
    b1123 := true;
    b1124 := true;
    b1125 := true;
    b1126 := true;
    b1127 := true;
    b1128 := true;
    b1129 := true;
    b1130 := true;
    b1131 := true;
    b1132 := true;
    b1133 := true;
    b1134 := true;
    b1135 := true;
    b1136 := true;
    b1137 := true;
    b1138 := true;
    b1139 := true;
    b1140 := true;
    b1141 := true;
    b1142 := true;
    b1143 := true;
    b1144 := true;
    b1145 := true;
    b1146 := true;
    b1147 := true;
    b1148 := true;
    b1149 := (b1084 AND (b1117 AND (b1118 AND (b1119 AND (b1120 AND (b1121 AND (b1122 AND (b1123 AND (b1124 AND (b1125 AND (b1126 AND (b1127 AND (b1128 AND (b1129 AND (b1130 AND (b1131 AND (b1132 AND (b1133 AND (b1134 AND (b1135 AND (b1136 AND (b1137 AND (b1138 AND (b1139 AND (b1140 AND (b1141 AND (b1142 AND (b1143 AND (b1144 AND (b1145 AND (b1146 AND (b1147 AND b1148))))))))))))))))))))))))))))))));
    null;
    null;
    r1151 := "0";
    null;
    r1152 := (r1151);
    r1153 := "0";
    null;
    r1154 := (r1153);
    r1155 := "0";
    null;
    r1156 := (r1155);
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    r1150 := (r1152 & r1154 & r1156 & r1085 & r1086 & r1087 & r1088 & r1089 & r1090 & r1091 & r1092 & r1093 & r1094 & r1095 & r1096 & r1097 & r1098 & r1099 & r1100 & r1101 & r1102 & r1103 & r1104 & r1105 & r1106 & r1107 & r1108 & r1109 & r1110 & r1111 & r1112 & r1113);
    r1083 := r1150;
    return r1083;
  end rewire_RWPrelude.shiftR3_1081;
  function rewire_RWPrelude.rotateR18_1009(r1010 : std_logic_vector) return std_logic_vector
  is
    variable r1078 : std_logic_vector(0 to 31) := (others => '0');
    variable b1077 : boolean := false;
    variable b1076 : boolean := false;
    variable b1075 : boolean := false;
    variable b1074 : boolean := false;
    variable b1073 : boolean := false;
    variable b1072 : boolean := false;
    variable b1071 : boolean := false;
    variable b1070 : boolean := false;
    variable b1069 : boolean := false;
    variable b1068 : boolean := false;
    variable b1067 : boolean := false;
    variable b1066 : boolean := false;
    variable b1065 : boolean := false;
    variable b1064 : boolean := false;
    variable b1063 : boolean := false;
    variable b1062 : boolean := false;
    variable b1061 : boolean := false;
    variable b1060 : boolean := false;
    variable b1059 : boolean := false;
    variable b1058 : boolean := false;
    variable b1057 : boolean := false;
    variable b1056 : boolean := false;
    variable b1055 : boolean := false;
    variable b1054 : boolean := false;
    variable b1053 : boolean := false;
    variable b1052 : boolean := false;
    variable b1051 : boolean := false;
    variable b1050 : boolean := false;
    variable b1049 : boolean := false;
    variable b1048 : boolean := false;
    variable b1047 : boolean := false;
    variable b1046 : boolean := false;
    variable b1045 : boolean := false;
    variable r1044 : std_logic_vector(0 to 0) := (others => '0');
    variable r1043 : std_logic_vector(0 to 0) := (others => '0');
    variable r1042 : std_logic_vector(0 to 0) := (others => '0');
    variable r1041 : std_logic_vector(0 to 0) := (others => '0');
    variable r1040 : std_logic_vector(0 to 0) := (others => '0');
    variable r1039 : std_logic_vector(0 to 0) := (others => '0');
    variable r1038 : std_logic_vector(0 to 0) := (others => '0');
    variable r1037 : std_logic_vector(0 to 0) := (others => '0');
    variable r1036 : std_logic_vector(0 to 0) := (others => '0');
    variable r1035 : std_logic_vector(0 to 0) := (others => '0');
    variable r1034 : std_logic_vector(0 to 0) := (others => '0');
    variable r1033 : std_logic_vector(0 to 0) := (others => '0');
    variable r1032 : std_logic_vector(0 to 0) := (others => '0');
    variable r1031 : std_logic_vector(0 to 0) := (others => '0');
    variable r1030 : std_logic_vector(0 to 0) := (others => '0');
    variable r1029 : std_logic_vector(0 to 0) := (others => '0');
    variable r1028 : std_logic_vector(0 to 0) := (others => '0');
    variable r1027 : std_logic_vector(0 to 0) := (others => '0');
    variable r1026 : std_logic_vector(0 to 0) := (others => '0');
    variable r1025 : std_logic_vector(0 to 0) := (others => '0');
    variable r1024 : std_logic_vector(0 to 0) := (others => '0');
    variable r1023 : std_logic_vector(0 to 0) := (others => '0');
    variable r1022 : std_logic_vector(0 to 0) := (others => '0');
    variable r1021 : std_logic_vector(0 to 0) := (others => '0');
    variable r1020 : std_logic_vector(0 to 0) := (others => '0');
    variable r1019 : std_logic_vector(0 to 0) := (others => '0');
    variable r1018 : std_logic_vector(0 to 0) := (others => '0');
    variable r1017 : std_logic_vector(0 to 0) := (others => '0');
    variable r1016 : std_logic_vector(0 to 0) := (others => '0');
    variable r1015 : std_logic_vector(0 to 0) := (others => '0');
    variable r1014 : std_logic_vector(0 to 0) := (others => '0');
    variable r1013 : std_logic_vector(0 to 0) := (others => '0');
    variable b1012 : boolean := false;
    variable r1011 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    b1012 := true;
    r1013 := r1010(0 to 0);
    r1014 := r1010(1 to 1);
    r1015 := r1010(2 to 2);
    r1016 := r1010(3 to 3);
    r1017 := r1010(4 to 4);
    r1018 := r1010(5 to 5);
    r1019 := r1010(6 to 6);
    r1020 := r1010(7 to 7);
    r1021 := r1010(8 to 8);
    r1022 := r1010(9 to 9);
    r1023 := r1010(10 to 10);
    r1024 := r1010(11 to 11);
    r1025 := r1010(12 to 12);
    r1026 := r1010(13 to 13);
    r1027 := r1010(14 to 14);
    r1028 := r1010(15 to 15);
    r1029 := r1010(16 to 16);
    r1030 := r1010(17 to 17);
    r1031 := r1010(18 to 18);
    r1032 := r1010(19 to 19);
    r1033 := r1010(20 to 20);
    r1034 := r1010(21 to 21);
    r1035 := r1010(22 to 22);
    r1036 := r1010(23 to 23);
    r1037 := r1010(24 to 24);
    r1038 := r1010(25 to 25);
    r1039 := r1010(26 to 26);
    r1040 := r1010(27 to 27);
    r1041 := r1010(28 to 28);
    r1042 := r1010(29 to 29);
    r1043 := r1010(30 to 30);
    r1044 := r1010(31 to 31);
    b1045 := true;
    b1046 := true;
    b1047 := true;
    b1048 := true;
    b1049 := true;
    b1050 := true;
    b1051 := true;
    b1052 := true;
    b1053 := true;
    b1054 := true;
    b1055 := true;
    b1056 := true;
    b1057 := true;
    b1058 := true;
    b1059 := true;
    b1060 := true;
    b1061 := true;
    b1062 := true;
    b1063 := true;
    b1064 := true;
    b1065 := true;
    b1066 := true;
    b1067 := true;
    b1068 := true;
    b1069 := true;
    b1070 := true;
    b1071 := true;
    b1072 := true;
    b1073 := true;
    b1074 := true;
    b1075 := true;
    b1076 := true;
    b1077 := (b1012 AND (b1045 AND (b1046 AND (b1047 AND (b1048 AND (b1049 AND (b1050 AND (b1051 AND (b1052 AND (b1053 AND (b1054 AND (b1055 AND (b1056 AND (b1057 AND (b1058 AND (b1059 AND (b1060 AND (b1061 AND (b1062 AND (b1063 AND (b1064 AND (b1065 AND (b1066 AND (b1067 AND (b1068 AND (b1069 AND (b1070 AND (b1071 AND (b1072 AND (b1073 AND (b1074 AND (b1075 AND b1076))))))))))))))))))))))))))))))));
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    r1078 := (r1027 & r1028 & r1029 & r1030 & r1031 & r1032 & r1033 & r1034 & r1035 & r1036 & r1037 & r1038 & r1039 & r1040 & r1041 & r1042 & r1043 & r1044 & r1013 & r1014 & r1015 & r1016 & r1017 & r1018 & r1019 & r1020 & r1021 & r1022 & r1023 & r1024 & r1025 & r1026);
    r1011 := r1078;
    return r1011;
  end rewire_RWPrelude.rotateR18_1009;
  function rewire_RWPrelude.rotateR7_938(r939 : std_logic_vector) return std_logic_vector
  is
    variable r1007 : std_logic_vector(0 to 31) := (others => '0');
    variable b1006 : boolean := false;
    variable b1005 : boolean := false;
    variable b1004 : boolean := false;
    variable b1003 : boolean := false;
    variable b1002 : boolean := false;
    variable b1001 : boolean := false;
    variable b1000 : boolean := false;
    variable b999 : boolean := false;
    variable b998 : boolean := false;
    variable b997 : boolean := false;
    variable b996 : boolean := false;
    variable b995 : boolean := false;
    variable b994 : boolean := false;
    variable b993 : boolean := false;
    variable b992 : boolean := false;
    variable b991 : boolean := false;
    variable b990 : boolean := false;
    variable b989 : boolean := false;
    variable b988 : boolean := false;
    variable b987 : boolean := false;
    variable b986 : boolean := false;
    variable b985 : boolean := false;
    variable b984 : boolean := false;
    variable b983 : boolean := false;
    variable b982 : boolean := false;
    variable b981 : boolean := false;
    variable b980 : boolean := false;
    variable b979 : boolean := false;
    variable b978 : boolean := false;
    variable b977 : boolean := false;
    variable b976 : boolean := false;
    variable b975 : boolean := false;
    variable b974 : boolean := false;
    variable r973 : std_logic_vector(0 to 0) := (others => '0');
    variable r972 : std_logic_vector(0 to 0) := (others => '0');
    variable r971 : std_logic_vector(0 to 0) := (others => '0');
    variable r970 : std_logic_vector(0 to 0) := (others => '0');
    variable r969 : std_logic_vector(0 to 0) := (others => '0');
    variable r968 : std_logic_vector(0 to 0) := (others => '0');
    variable r967 : std_logic_vector(0 to 0) := (others => '0');
    variable r966 : std_logic_vector(0 to 0) := (others => '0');
    variable r965 : std_logic_vector(0 to 0) := (others => '0');
    variable r964 : std_logic_vector(0 to 0) := (others => '0');
    variable r963 : std_logic_vector(0 to 0) := (others => '0');
    variable r962 : std_logic_vector(0 to 0) := (others => '0');
    variable r961 : std_logic_vector(0 to 0) := (others => '0');
    variable r960 : std_logic_vector(0 to 0) := (others => '0');
    variable r959 : std_logic_vector(0 to 0) := (others => '0');
    variable r958 : std_logic_vector(0 to 0) := (others => '0');
    variable r957 : std_logic_vector(0 to 0) := (others => '0');
    variable r956 : std_logic_vector(0 to 0) := (others => '0');
    variable r955 : std_logic_vector(0 to 0) := (others => '0');
    variable r954 : std_logic_vector(0 to 0) := (others => '0');
    variable r953 : std_logic_vector(0 to 0) := (others => '0');
    variable r952 : std_logic_vector(0 to 0) := (others => '0');
    variable r951 : std_logic_vector(0 to 0) := (others => '0');
    variable r950 : std_logic_vector(0 to 0) := (others => '0');
    variable r949 : std_logic_vector(0 to 0) := (others => '0');
    variable r948 : std_logic_vector(0 to 0) := (others => '0');
    variable r947 : std_logic_vector(0 to 0) := (others => '0');
    variable r946 : std_logic_vector(0 to 0) := (others => '0');
    variable r945 : std_logic_vector(0 to 0) := (others => '0');
    variable r944 : std_logic_vector(0 to 0) := (others => '0');
    variable r943 : std_logic_vector(0 to 0) := (others => '0');
    variable r942 : std_logic_vector(0 to 0) := (others => '0');
    variable b941 : boolean := false;
    variable r940 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    b941 := true;
    r942 := r939(0 to 0);
    r943 := r939(1 to 1);
    r944 := r939(2 to 2);
    r945 := r939(3 to 3);
    r946 := r939(4 to 4);
    r947 := r939(5 to 5);
    r948 := r939(6 to 6);
    r949 := r939(7 to 7);
    r950 := r939(8 to 8);
    r951 := r939(9 to 9);
    r952 := r939(10 to 10);
    r953 := r939(11 to 11);
    r954 := r939(12 to 12);
    r955 := r939(13 to 13);
    r956 := r939(14 to 14);
    r957 := r939(15 to 15);
    r958 := r939(16 to 16);
    r959 := r939(17 to 17);
    r960 := r939(18 to 18);
    r961 := r939(19 to 19);
    r962 := r939(20 to 20);
    r963 := r939(21 to 21);
    r964 := r939(22 to 22);
    r965 := r939(23 to 23);
    r966 := r939(24 to 24);
    r967 := r939(25 to 25);
    r968 := r939(26 to 26);
    r969 := r939(27 to 27);
    r970 := r939(28 to 28);
    r971 := r939(29 to 29);
    r972 := r939(30 to 30);
    r973 := r939(31 to 31);
    b974 := true;
    b975 := true;
    b976 := true;
    b977 := true;
    b978 := true;
    b979 := true;
    b980 := true;
    b981 := true;
    b982 := true;
    b983 := true;
    b984 := true;
    b985 := true;
    b986 := true;
    b987 := true;
    b988 := true;
    b989 := true;
    b990 := true;
    b991 := true;
    b992 := true;
    b993 := true;
    b994 := true;
    b995 := true;
    b996 := true;
    b997 := true;
    b998 := true;
    b999 := true;
    b1000 := true;
    b1001 := true;
    b1002 := true;
    b1003 := true;
    b1004 := true;
    b1005 := true;
    b1006 := (b941 AND (b974 AND (b975 AND (b976 AND (b977 AND (b978 AND (b979 AND (b980 AND (b981 AND (b982 AND (b983 AND (b984 AND (b985 AND (b986 AND (b987 AND (b988 AND (b989 AND (b990 AND (b991 AND (b992 AND (b993 AND (b994 AND (b995 AND (b996 AND (b997 AND (b998 AND (b999 AND (b1000 AND (b1001 AND (b1002 AND (b1003 AND (b1004 AND b1005))))))))))))))))))))))))))))))));
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    r1007 := (r967 & r968 & r969 & r970 & r971 & r972 & r973 & r942 & r943 & r944 & r945 & r946 & r947 & r948 & r949 & r950 & r951 & r952 & r953 & r954 & r955 & r956 & r957 & r958 & r959 & r960 & r961 & r962 & r963 & r964 & r965 & r966);
    r940 := r1007;
    return r940;
  end rewire_RWPrelude.rotateR7_938;
  function rewire_Main.sigma1_697(r698 : std_logic_vector) return std_logic_vector
  is
    variable r933 : std_logic_vector(0 to 31) := (others => '0');
    variable r932 : std_logic_vector(0 to 31) := (others => '0');
    variable r843 : std_logic_vector(0 to 31) := (others => '0');
    variable r841 : std_logic_vector(0 to 31) := (others => '0');
    variable r840 : std_logic_vector(0 to 31) := (others => '0');
    variable r771 : std_logic_vector(0 to 31) := (others => '0');
    variable r769 : std_logic_vector(0 to 31) := (others => '0');
    variable r700 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    r769 := rewire_RWPrelude.rotateR17_699(r698);
    null;
    r840 := rewire_RWPrelude.rotateR19_770(r698);
    r841 := w32Xor(r769,r840);
    null;
    r932 := rewire_RWPrelude.shiftR10_842(r698);
    r933 := w32Xor(r841,r932);
    return r933;
  end rewire_Main.sigma1_697;
  function rewire_RWPrelude.shiftR10_842(r843 : std_logic_vector) return std_logic_vector
  is
    variable r931 : std_logic_vector(0 to 0) := (others => '0');
    variable r930 : std_logic_vector(0 to 0) := (others => '0');
    variable r929 : std_logic_vector(0 to 0) := (others => '0');
    variable r928 : std_logic_vector(0 to 0) := (others => '0');
    variable r927 : std_logic_vector(0 to 0) := (others => '0');
    variable r926 : std_logic_vector(0 to 0) := (others => '0');
    variable r925 : std_logic_vector(0 to 0) := (others => '0');
    variable r924 : std_logic_vector(0 to 0) := (others => '0');
    variable r923 : std_logic_vector(0 to 0) := (others => '0');
    variable r922 : std_logic_vector(0 to 0) := (others => '0');
    variable r921 : std_logic_vector(0 to 0) := (others => '0');
    variable r920 : std_logic_vector(0 to 0) := (others => '0');
    variable r919 : std_logic_vector(0 to 0) := (others => '0');
    variable r918 : std_logic_vector(0 to 0) := (others => '0');
    variable r917 : std_logic_vector(0 to 0) := (others => '0');
    variable r916 : std_logic_vector(0 to 0) := (others => '0');
    variable r915 : std_logic_vector(0 to 0) := (others => '0');
    variable r914 : std_logic_vector(0 to 0) := (others => '0');
    variable r913 : std_logic_vector(0 to 0) := (others => '0');
    variable r912 : std_logic_vector(0 to 0) := (others => '0');
    variable r911 : std_logic_vector(0 to 31) := (others => '0');
    variable b910 : boolean := false;
    variable b909 : boolean := false;
    variable b908 : boolean := false;
    variable b907 : boolean := false;
    variable b906 : boolean := false;
    variable b905 : boolean := false;
    variable b904 : boolean := false;
    variable b903 : boolean := false;
    variable b902 : boolean := false;
    variable b901 : boolean := false;
    variable b900 : boolean := false;
    variable b899 : boolean := false;
    variable b898 : boolean := false;
    variable b897 : boolean := false;
    variable b896 : boolean := false;
    variable b895 : boolean := false;
    variable b894 : boolean := false;
    variable b893 : boolean := false;
    variable b892 : boolean := false;
    variable b891 : boolean := false;
    variable b890 : boolean := false;
    variable b889 : boolean := false;
    variable b888 : boolean := false;
    variable b887 : boolean := false;
    variable b886 : boolean := false;
    variable b885 : boolean := false;
    variable b884 : boolean := false;
    variable b883 : boolean := false;
    variable b882 : boolean := false;
    variable b881 : boolean := false;
    variable b880 : boolean := false;
    variable b879 : boolean := false;
    variable b878 : boolean := false;
    variable r877 : std_logic_vector(0 to 0) := (others => '0');
    variable r876 : std_logic_vector(0 to 0) := (others => '0');
    variable r875 : std_logic_vector(0 to 0) := (others => '0');
    variable r874 : std_logic_vector(0 to 0) := (others => '0');
    variable r873 : std_logic_vector(0 to 0) := (others => '0');
    variable r872 : std_logic_vector(0 to 0) := (others => '0');
    variable r871 : std_logic_vector(0 to 0) := (others => '0');
    variable r870 : std_logic_vector(0 to 0) := (others => '0');
    variable r869 : std_logic_vector(0 to 0) := (others => '0');
    variable r868 : std_logic_vector(0 to 0) := (others => '0');
    variable r867 : std_logic_vector(0 to 0) := (others => '0');
    variable r866 : std_logic_vector(0 to 0) := (others => '0');
    variable r865 : std_logic_vector(0 to 0) := (others => '0');
    variable r864 : std_logic_vector(0 to 0) := (others => '0');
    variable r863 : std_logic_vector(0 to 0) := (others => '0');
    variable r862 : std_logic_vector(0 to 0) := (others => '0');
    variable r861 : std_logic_vector(0 to 0) := (others => '0');
    variable r860 : std_logic_vector(0 to 0) := (others => '0');
    variable r859 : std_logic_vector(0 to 0) := (others => '0');
    variable r858 : std_logic_vector(0 to 0) := (others => '0');
    variable r857 : std_logic_vector(0 to 0) := (others => '0');
    variable r856 : std_logic_vector(0 to 0) := (others => '0');
    variable r855 : std_logic_vector(0 to 0) := (others => '0');
    variable r854 : std_logic_vector(0 to 0) := (others => '0');
    variable r853 : std_logic_vector(0 to 0) := (others => '0');
    variable r852 : std_logic_vector(0 to 0) := (others => '0');
    variable r851 : std_logic_vector(0 to 0) := (others => '0');
    variable r850 : std_logic_vector(0 to 0) := (others => '0');
    variable r849 : std_logic_vector(0 to 0) := (others => '0');
    variable r848 : std_logic_vector(0 to 0) := (others => '0');
    variable r847 : std_logic_vector(0 to 0) := (others => '0');
    variable r846 : std_logic_vector(0 to 0) := (others => '0');
    variable b845 : boolean := false;
    variable r844 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    b845 := true;
    r846 := r843(0 to 0);
    r847 := r843(1 to 1);
    r848 := r843(2 to 2);
    r849 := r843(3 to 3);
    r850 := r843(4 to 4);
    r851 := r843(5 to 5);
    r852 := r843(6 to 6);
    r853 := r843(7 to 7);
    r854 := r843(8 to 8);
    r855 := r843(9 to 9);
    r856 := r843(10 to 10);
    r857 := r843(11 to 11);
    r858 := r843(12 to 12);
    r859 := r843(13 to 13);
    r860 := r843(14 to 14);
    r861 := r843(15 to 15);
    r862 := r843(16 to 16);
    r863 := r843(17 to 17);
    r864 := r843(18 to 18);
    r865 := r843(19 to 19);
    r866 := r843(20 to 20);
    r867 := r843(21 to 21);
    r868 := r843(22 to 22);
    r869 := r843(23 to 23);
    r870 := r843(24 to 24);
    r871 := r843(25 to 25);
    r872 := r843(26 to 26);
    r873 := r843(27 to 27);
    r874 := r843(28 to 28);
    r875 := r843(29 to 29);
    r876 := r843(30 to 30);
    r877 := r843(31 to 31);
    b878 := true;
    b879 := true;
    b880 := true;
    b881 := true;
    b882 := true;
    b883 := true;
    b884 := true;
    b885 := true;
    b886 := true;
    b887 := true;
    b888 := true;
    b889 := true;
    b890 := true;
    b891 := true;
    b892 := true;
    b893 := true;
    b894 := true;
    b895 := true;
    b896 := true;
    b897 := true;
    b898 := true;
    b899 := true;
    b900 := true;
    b901 := true;
    b902 := true;
    b903 := true;
    b904 := true;
    b905 := true;
    b906 := true;
    b907 := true;
    b908 := true;
    b909 := true;
    b910 := (b845 AND (b878 AND (b879 AND (b880 AND (b881 AND (b882 AND (b883 AND (b884 AND (b885 AND (b886 AND (b887 AND (b888 AND (b889 AND (b890 AND (b891 AND (b892 AND (b893 AND (b894 AND (b895 AND (b896 AND (b897 AND (b898 AND (b899 AND (b900 AND (b901 AND (b902 AND (b903 AND (b904 AND (b905 AND (b906 AND (b907 AND (b908 AND b909))))))))))))))))))))))))))))))));
    null;
    null;
    r912 := "0";
    null;
    r913 := (r912);
    r914 := "0";
    null;
    r915 := (r914);
    r916 := "0";
    null;
    r917 := (r916);
    r918 := "0";
    null;
    r919 := (r918);
    r920 := "0";
    null;
    r921 := (r920);
    r922 := "0";
    null;
    r923 := (r922);
    r924 := "0";
    null;
    r925 := (r924);
    r926 := "0";
    null;
    r927 := (r926);
    r928 := "0";
    null;
    r929 := (r928);
    r930 := "0";
    null;
    r931 := (r930);
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    r911 := (r913 & r915 & r917 & r919 & r921 & r923 & r925 & r927 & r929 & r931 & r846 & r847 & r848 & r849 & r850 & r851 & r852 & r853 & r854 & r855 & r856 & r857 & r858 & r859 & r860 & r861 & r862 & r863 & r864 & r865 & r866 & r867);
    r844 := r911;
    return r844;
  end rewire_RWPrelude.shiftR10_842;
  function rewire_RWPrelude.rotateR19_770(r771 : std_logic_vector) return std_logic_vector
  is
    variable r839 : std_logic_vector(0 to 31) := (others => '0');
    variable b838 : boolean := false;
    variable b837 : boolean := false;
    variable b836 : boolean := false;
    variable b835 : boolean := false;
    variable b834 : boolean := false;
    variable b833 : boolean := false;
    variable b832 : boolean := false;
    variable b831 : boolean := false;
    variable b830 : boolean := false;
    variable b829 : boolean := false;
    variable b828 : boolean := false;
    variable b827 : boolean := false;
    variable b826 : boolean := false;
    variable b825 : boolean := false;
    variable b824 : boolean := false;
    variable b823 : boolean := false;
    variable b822 : boolean := false;
    variable b821 : boolean := false;
    variable b820 : boolean := false;
    variable b819 : boolean := false;
    variable b818 : boolean := false;
    variable b817 : boolean := false;
    variable b816 : boolean := false;
    variable b815 : boolean := false;
    variable b814 : boolean := false;
    variable b813 : boolean := false;
    variable b812 : boolean := false;
    variable b811 : boolean := false;
    variable b810 : boolean := false;
    variable b809 : boolean := false;
    variable b808 : boolean := false;
    variable b807 : boolean := false;
    variable b806 : boolean := false;
    variable r805 : std_logic_vector(0 to 0) := (others => '0');
    variable r804 : std_logic_vector(0 to 0) := (others => '0');
    variable r803 : std_logic_vector(0 to 0) := (others => '0');
    variable r802 : std_logic_vector(0 to 0) := (others => '0');
    variable r801 : std_logic_vector(0 to 0) := (others => '0');
    variable r800 : std_logic_vector(0 to 0) := (others => '0');
    variable r799 : std_logic_vector(0 to 0) := (others => '0');
    variable r798 : std_logic_vector(0 to 0) := (others => '0');
    variable r797 : std_logic_vector(0 to 0) := (others => '0');
    variable r796 : std_logic_vector(0 to 0) := (others => '0');
    variable r795 : std_logic_vector(0 to 0) := (others => '0');
    variable r794 : std_logic_vector(0 to 0) := (others => '0');
    variable r793 : std_logic_vector(0 to 0) := (others => '0');
    variable r792 : std_logic_vector(0 to 0) := (others => '0');
    variable r791 : std_logic_vector(0 to 0) := (others => '0');
    variable r790 : std_logic_vector(0 to 0) := (others => '0');
    variable r789 : std_logic_vector(0 to 0) := (others => '0');
    variable r788 : std_logic_vector(0 to 0) := (others => '0');
    variable r787 : std_logic_vector(0 to 0) := (others => '0');
    variable r786 : std_logic_vector(0 to 0) := (others => '0');
    variable r785 : std_logic_vector(0 to 0) := (others => '0');
    variable r784 : std_logic_vector(0 to 0) := (others => '0');
    variable r783 : std_logic_vector(0 to 0) := (others => '0');
    variable r782 : std_logic_vector(0 to 0) := (others => '0');
    variable r781 : std_logic_vector(0 to 0) := (others => '0');
    variable r780 : std_logic_vector(0 to 0) := (others => '0');
    variable r779 : std_logic_vector(0 to 0) := (others => '0');
    variable r778 : std_logic_vector(0 to 0) := (others => '0');
    variable r777 : std_logic_vector(0 to 0) := (others => '0');
    variable r776 : std_logic_vector(0 to 0) := (others => '0');
    variable r775 : std_logic_vector(0 to 0) := (others => '0');
    variable r774 : std_logic_vector(0 to 0) := (others => '0');
    variable b773 : boolean := false;
    variable r772 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    b773 := true;
    r774 := r771(0 to 0);
    r775 := r771(1 to 1);
    r776 := r771(2 to 2);
    r777 := r771(3 to 3);
    r778 := r771(4 to 4);
    r779 := r771(5 to 5);
    r780 := r771(6 to 6);
    r781 := r771(7 to 7);
    r782 := r771(8 to 8);
    r783 := r771(9 to 9);
    r784 := r771(10 to 10);
    r785 := r771(11 to 11);
    r786 := r771(12 to 12);
    r787 := r771(13 to 13);
    r788 := r771(14 to 14);
    r789 := r771(15 to 15);
    r790 := r771(16 to 16);
    r791 := r771(17 to 17);
    r792 := r771(18 to 18);
    r793 := r771(19 to 19);
    r794 := r771(20 to 20);
    r795 := r771(21 to 21);
    r796 := r771(22 to 22);
    r797 := r771(23 to 23);
    r798 := r771(24 to 24);
    r799 := r771(25 to 25);
    r800 := r771(26 to 26);
    r801 := r771(27 to 27);
    r802 := r771(28 to 28);
    r803 := r771(29 to 29);
    r804 := r771(30 to 30);
    r805 := r771(31 to 31);
    b806 := true;
    b807 := true;
    b808 := true;
    b809 := true;
    b810 := true;
    b811 := true;
    b812 := true;
    b813 := true;
    b814 := true;
    b815 := true;
    b816 := true;
    b817 := true;
    b818 := true;
    b819 := true;
    b820 := true;
    b821 := true;
    b822 := true;
    b823 := true;
    b824 := true;
    b825 := true;
    b826 := true;
    b827 := true;
    b828 := true;
    b829 := true;
    b830 := true;
    b831 := true;
    b832 := true;
    b833 := true;
    b834 := true;
    b835 := true;
    b836 := true;
    b837 := true;
    b838 := (b773 AND (b806 AND (b807 AND (b808 AND (b809 AND (b810 AND (b811 AND (b812 AND (b813 AND (b814 AND (b815 AND (b816 AND (b817 AND (b818 AND (b819 AND (b820 AND (b821 AND (b822 AND (b823 AND (b824 AND (b825 AND (b826 AND (b827 AND (b828 AND (b829 AND (b830 AND (b831 AND (b832 AND (b833 AND (b834 AND (b835 AND (b836 AND b837))))))))))))))))))))))))))))))));
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    r839 := (r787 & r788 & r789 & r790 & r791 & r792 & r793 & r794 & r795 & r796 & r797 & r798 & r799 & r800 & r801 & r802 & r803 & r804 & r805 & r774 & r775 & r776 & r777 & r778 & r779 & r780 & r781 & r782 & r783 & r784 & r785 & r786);
    r772 := r839;
    return r772;
  end rewire_RWPrelude.rotateR19_770;
  function rewire_RWPrelude.rotateR17_699(r700 : std_logic_vector) return std_logic_vector
  is
    variable r768 : std_logic_vector(0 to 31) := (others => '0');
    variable b767 : boolean := false;
    variable b766 : boolean := false;
    variable b765 : boolean := false;
    variable b764 : boolean := false;
    variable b763 : boolean := false;
    variable b762 : boolean := false;
    variable b761 : boolean := false;
    variable b760 : boolean := false;
    variable b759 : boolean := false;
    variable b758 : boolean := false;
    variable b757 : boolean := false;
    variable b756 : boolean := false;
    variable b755 : boolean := false;
    variable b754 : boolean := false;
    variable b753 : boolean := false;
    variable b752 : boolean := false;
    variable b751 : boolean := false;
    variable b750 : boolean := false;
    variable b749 : boolean := false;
    variable b748 : boolean := false;
    variable b747 : boolean := false;
    variable b746 : boolean := false;
    variable b745 : boolean := false;
    variable b744 : boolean := false;
    variable b743 : boolean := false;
    variable b742 : boolean := false;
    variable b741 : boolean := false;
    variable b740 : boolean := false;
    variable b739 : boolean := false;
    variable b738 : boolean := false;
    variable b737 : boolean := false;
    variable b736 : boolean := false;
    variable b735 : boolean := false;
    variable r734 : std_logic_vector(0 to 0) := (others => '0');
    variable r733 : std_logic_vector(0 to 0) := (others => '0');
    variable r732 : std_logic_vector(0 to 0) := (others => '0');
    variable r731 : std_logic_vector(0 to 0) := (others => '0');
    variable r730 : std_logic_vector(0 to 0) := (others => '0');
    variable r729 : std_logic_vector(0 to 0) := (others => '0');
    variable r728 : std_logic_vector(0 to 0) := (others => '0');
    variable r727 : std_logic_vector(0 to 0) := (others => '0');
    variable r726 : std_logic_vector(0 to 0) := (others => '0');
    variable r725 : std_logic_vector(0 to 0) := (others => '0');
    variable r724 : std_logic_vector(0 to 0) := (others => '0');
    variable r723 : std_logic_vector(0 to 0) := (others => '0');
    variable r722 : std_logic_vector(0 to 0) := (others => '0');
    variable r721 : std_logic_vector(0 to 0) := (others => '0');
    variable r720 : std_logic_vector(0 to 0) := (others => '0');
    variable r719 : std_logic_vector(0 to 0) := (others => '0');
    variable r718 : std_logic_vector(0 to 0) := (others => '0');
    variable r717 : std_logic_vector(0 to 0) := (others => '0');
    variable r716 : std_logic_vector(0 to 0) := (others => '0');
    variable r715 : std_logic_vector(0 to 0) := (others => '0');
    variable r714 : std_logic_vector(0 to 0) := (others => '0');
    variable r713 : std_logic_vector(0 to 0) := (others => '0');
    variable r712 : std_logic_vector(0 to 0) := (others => '0');
    variable r711 : std_logic_vector(0 to 0) := (others => '0');
    variable r710 : std_logic_vector(0 to 0) := (others => '0');
    variable r709 : std_logic_vector(0 to 0) := (others => '0');
    variable r708 : std_logic_vector(0 to 0) := (others => '0');
    variable r707 : std_logic_vector(0 to 0) := (others => '0');
    variable r706 : std_logic_vector(0 to 0) := (others => '0');
    variable r705 : std_logic_vector(0 to 0) := (others => '0');
    variable r704 : std_logic_vector(0 to 0) := (others => '0');
    variable r703 : std_logic_vector(0 to 0) := (others => '0');
    variable b702 : boolean := false;
    variable r701 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    b702 := true;
    r703 := r700(0 to 0);
    r704 := r700(1 to 1);
    r705 := r700(2 to 2);
    r706 := r700(3 to 3);
    r707 := r700(4 to 4);
    r708 := r700(5 to 5);
    r709 := r700(6 to 6);
    r710 := r700(7 to 7);
    r711 := r700(8 to 8);
    r712 := r700(9 to 9);
    r713 := r700(10 to 10);
    r714 := r700(11 to 11);
    r715 := r700(12 to 12);
    r716 := r700(13 to 13);
    r717 := r700(14 to 14);
    r718 := r700(15 to 15);
    r719 := r700(16 to 16);
    r720 := r700(17 to 17);
    r721 := r700(18 to 18);
    r722 := r700(19 to 19);
    r723 := r700(20 to 20);
    r724 := r700(21 to 21);
    r725 := r700(22 to 22);
    r726 := r700(23 to 23);
    r727 := r700(24 to 24);
    r728 := r700(25 to 25);
    r729 := r700(26 to 26);
    r730 := r700(27 to 27);
    r731 := r700(28 to 28);
    r732 := r700(29 to 29);
    r733 := r700(30 to 30);
    r734 := r700(31 to 31);
    b735 := true;
    b736 := true;
    b737 := true;
    b738 := true;
    b739 := true;
    b740 := true;
    b741 := true;
    b742 := true;
    b743 := true;
    b744 := true;
    b745 := true;
    b746 := true;
    b747 := true;
    b748 := true;
    b749 := true;
    b750 := true;
    b751 := true;
    b752 := true;
    b753 := true;
    b754 := true;
    b755 := true;
    b756 := true;
    b757 := true;
    b758 := true;
    b759 := true;
    b760 := true;
    b761 := true;
    b762 := true;
    b763 := true;
    b764 := true;
    b765 := true;
    b766 := true;
    b767 := (b702 AND (b735 AND (b736 AND (b737 AND (b738 AND (b739 AND (b740 AND (b741 AND (b742 AND (b743 AND (b744 AND (b745 AND (b746 AND (b747 AND (b748 AND (b749 AND (b750 AND (b751 AND (b752 AND (b753 AND (b754 AND (b755 AND (b756 AND (b757 AND (b758 AND (b759 AND (b760 AND (b761 AND (b762 AND (b763 AND (b764 AND (b765 AND b766))))))))))))))))))))))))))))))));
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    null;
    r768 := (r718 & r719 & r720 & r721 & r722 & r723 & r724 & r725 & r726 & r727 & r728 & r729 & r730 & r731 & r732 & r733 & r734 & r703 & r704 & r705 & r706 & r707 & r708 & r709 & r710 & r711 & r712 & r713 & r714 & r715 & r716 & r717);
    r701 := r768;
    return r701;
  end rewire_RWPrelude.rotateR17_699;
  function rewire_Main.initialSHA256State_24 return std_logic_vector
  is
    variable r561 : std_logic_vector(0 to 31) := (others => '0');
    variable r494 : std_logic_vector(0 to 31) := (others => '0');
    variable r427 : std_logic_vector(0 to 31) := (others => '0');
    variable r360 : std_logic_vector(0 to 31) := (others => '0');
    variable r293 : std_logic_vector(0 to 31) := (others => '0');
    variable r226 : std_logic_vector(0 to 31) := (others => '0');
    variable r159 : std_logic_vector(0 to 31) := (others => '0');
    variable r92 : std_logic_vector(0 to 31) := (others => '0');
    variable r25 : std_logic_vector(0 to 255) := (others => '0');
  begin
    null;
    null;
    r92 := rewire_MetaprogrammingRW.w6a09e667_26;
    r159 := rewire_MetaprogrammingRW.wbb67ae85_93;
    r226 := rewire_MetaprogrammingRW.w3c6ef372_160;
    r293 := rewire_MetaprogrammingRW.wa54ff53a_227;
    r360 := rewire_MetaprogrammingRW.w510e527f_294;
    r427 := rewire_MetaprogrammingRW.w9b05688c_361;
    r494 := rewire_MetaprogrammingRW.w1f83d9ab_428;
    r561 := rewire_MetaprogrammingRW.w5be0cd19_495;
    r25 := (r92 & r159 & r226 & r293 & r360 & r427 & r494 & r561);
    return r25;
  end rewire_Main.initialSHA256State_24;
  function rewire_MetaprogrammingRW.w5be0cd19_495 return std_logic_vector
  is
    variable r560 : std_logic_vector(0 to 0) := (others => '0');
    variable r559 : std_logic_vector(0 to 0) := (others => '0');
    variable r558 : std_logic_vector(0 to 0) := (others => '0');
    variable r557 : std_logic_vector(0 to 0) := (others => '0');
    variable r556 : std_logic_vector(0 to 0) := (others => '0');
    variable r555 : std_logic_vector(0 to 0) := (others => '0');
    variable r554 : std_logic_vector(0 to 0) := (others => '0');
    variable r553 : std_logic_vector(0 to 0) := (others => '0');
    variable r552 : std_logic_vector(0 to 0) := (others => '0');
    variable r551 : std_logic_vector(0 to 0) := (others => '0');
    variable r550 : std_logic_vector(0 to 0) := (others => '0');
    variable r549 : std_logic_vector(0 to 0) := (others => '0');
    variable r548 : std_logic_vector(0 to 0) := (others => '0');
    variable r547 : std_logic_vector(0 to 0) := (others => '0');
    variable r546 : std_logic_vector(0 to 0) := (others => '0');
    variable r545 : std_logic_vector(0 to 0) := (others => '0');
    variable r544 : std_logic_vector(0 to 0) := (others => '0');
    variable r543 : std_logic_vector(0 to 0) := (others => '0');
    variable r542 : std_logic_vector(0 to 0) := (others => '0');
    variable r541 : std_logic_vector(0 to 0) := (others => '0');
    variable r540 : std_logic_vector(0 to 0) := (others => '0');
    variable r539 : std_logic_vector(0 to 0) := (others => '0');
    variable r538 : std_logic_vector(0 to 0) := (others => '0');
    variable r537 : std_logic_vector(0 to 0) := (others => '0');
    variable r536 : std_logic_vector(0 to 0) := (others => '0');
    variable r535 : std_logic_vector(0 to 0) := (others => '0');
    variable r534 : std_logic_vector(0 to 0) := (others => '0');
    variable r533 : std_logic_vector(0 to 0) := (others => '0');
    variable r532 : std_logic_vector(0 to 0) := (others => '0');
    variable r531 : std_logic_vector(0 to 0) := (others => '0');
    variable r530 : std_logic_vector(0 to 0) := (others => '0');
    variable r529 : std_logic_vector(0 to 0) := (others => '0');
    variable r528 : std_logic_vector(0 to 0) := (others => '0');
    variable r527 : std_logic_vector(0 to 0) := (others => '0');
    variable r526 : std_logic_vector(0 to 0) := (others => '0');
    variable r525 : std_logic_vector(0 to 0) := (others => '0');
    variable r524 : std_logic_vector(0 to 0) := (others => '0');
    variable r523 : std_logic_vector(0 to 0) := (others => '0');
    variable r522 : std_logic_vector(0 to 0) := (others => '0');
    variable r521 : std_logic_vector(0 to 0) := (others => '0');
    variable r520 : std_logic_vector(0 to 0) := (others => '0');
    variable r519 : std_logic_vector(0 to 0) := (others => '0');
    variable r518 : std_logic_vector(0 to 0) := (others => '0');
    variable r517 : std_logic_vector(0 to 0) := (others => '0');
    variable r516 : std_logic_vector(0 to 0) := (others => '0');
    variable r515 : std_logic_vector(0 to 0) := (others => '0');
    variable r514 : std_logic_vector(0 to 0) := (others => '0');
    variable r513 : std_logic_vector(0 to 0) := (others => '0');
    variable r512 : std_logic_vector(0 to 0) := (others => '0');
    variable r511 : std_logic_vector(0 to 0) := (others => '0');
    variable r510 : std_logic_vector(0 to 0) := (others => '0');
    variable r509 : std_logic_vector(0 to 0) := (others => '0');
    variable r508 : std_logic_vector(0 to 0) := (others => '0');
    variable r507 : std_logic_vector(0 to 0) := (others => '0');
    variable r506 : std_logic_vector(0 to 0) := (others => '0');
    variable r505 : std_logic_vector(0 to 0) := (others => '0');
    variable r504 : std_logic_vector(0 to 0) := (others => '0');
    variable r503 : std_logic_vector(0 to 0) := (others => '0');
    variable r502 : std_logic_vector(0 to 0) := (others => '0');
    variable r501 : std_logic_vector(0 to 0) := (others => '0');
    variable r500 : std_logic_vector(0 to 0) := (others => '0');
    variable r499 : std_logic_vector(0 to 0) := (others => '0');
    variable r498 : std_logic_vector(0 to 0) := (others => '0');
    variable r497 : std_logic_vector(0 to 0) := (others => '0');
    variable r496 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r497 := "0";
    null;
    r498 := (r497);
    r499 := "1";
    null;
    r500 := (r499);
    r501 := "0";
    null;
    r502 := (r501);
    r503 := "1";
    null;
    r504 := (r503);
    r505 := "1";
    null;
    r506 := (r505);
    r507 := "0";
    null;
    r508 := (r507);
    r509 := "1";
    null;
    r510 := (r509);
    r511 := "1";
    null;
    r512 := (r511);
    r513 := "1";
    null;
    r514 := (r513);
    r515 := "1";
    null;
    r516 := (r515);
    r517 := "1";
    null;
    r518 := (r517);
    r519 := "0";
    null;
    r520 := (r519);
    r521 := "0";
    null;
    r522 := (r521);
    r523 := "0";
    null;
    r524 := (r523);
    r525 := "0";
    null;
    r526 := (r525);
    r527 := "0";
    null;
    r528 := (r527);
    r529 := "1";
    null;
    r530 := (r529);
    r531 := "1";
    null;
    r532 := (r531);
    r533 := "0";
    null;
    r534 := (r533);
    r535 := "0";
    null;
    r536 := (r535);
    r537 := "1";
    null;
    r538 := (r537);
    r539 := "1";
    null;
    r540 := (r539);
    r541 := "0";
    null;
    r542 := (r541);
    r543 := "1";
    null;
    r544 := (r543);
    r545 := "0";
    null;
    r546 := (r545);
    r547 := "0";
    null;
    r548 := (r547);
    r549 := "0";
    null;
    r550 := (r549);
    r551 := "1";
    null;
    r552 := (r551);
    r553 := "1";
    null;
    r554 := (r553);
    r555 := "0";
    null;
    r556 := (r555);
    r557 := "0";
    null;
    r558 := (r557);
    r559 := "1";
    null;
    r560 := (r559);
    r496 := (r498 & r500 & r502 & r504 & r506 & r508 & r510 & r512 & r514 & r516 & r518 & r520 & r522 & r524 & r526 & r528 & r530 & r532 & r534 & r536 & r538 & r540 & r542 & r544 & r546 & r548 & r550 & r552 & r554 & r556 & r558 & r560);
    return r496;
  end rewire_MetaprogrammingRW.w5be0cd19_495;
  function rewire_MetaprogrammingRW.w1f83d9ab_428 return std_logic_vector
  is
    variable r493 : std_logic_vector(0 to 0) := (others => '0');
    variable r492 : std_logic_vector(0 to 0) := (others => '0');
    variable r491 : std_logic_vector(0 to 0) := (others => '0');
    variable r490 : std_logic_vector(0 to 0) := (others => '0');
    variable r489 : std_logic_vector(0 to 0) := (others => '0');
    variable r488 : std_logic_vector(0 to 0) := (others => '0');
    variable r487 : std_logic_vector(0 to 0) := (others => '0');
    variable r486 : std_logic_vector(0 to 0) := (others => '0');
    variable r485 : std_logic_vector(0 to 0) := (others => '0');
    variable r484 : std_logic_vector(0 to 0) := (others => '0');
    variable r483 : std_logic_vector(0 to 0) := (others => '0');
    variable r482 : std_logic_vector(0 to 0) := (others => '0');
    variable r481 : std_logic_vector(0 to 0) := (others => '0');
    variable r480 : std_logic_vector(0 to 0) := (others => '0');
    variable r479 : std_logic_vector(0 to 0) := (others => '0');
    variable r478 : std_logic_vector(0 to 0) := (others => '0');
    variable r477 : std_logic_vector(0 to 0) := (others => '0');
    variable r476 : std_logic_vector(0 to 0) := (others => '0');
    variable r475 : std_logic_vector(0 to 0) := (others => '0');
    variable r474 : std_logic_vector(0 to 0) := (others => '0');
    variable r473 : std_logic_vector(0 to 0) := (others => '0');
    variable r472 : std_logic_vector(0 to 0) := (others => '0');
    variable r471 : std_logic_vector(0 to 0) := (others => '0');
    variable r470 : std_logic_vector(0 to 0) := (others => '0');
    variable r469 : std_logic_vector(0 to 0) := (others => '0');
    variable r468 : std_logic_vector(0 to 0) := (others => '0');
    variable r467 : std_logic_vector(0 to 0) := (others => '0');
    variable r466 : std_logic_vector(0 to 0) := (others => '0');
    variable r465 : std_logic_vector(0 to 0) := (others => '0');
    variable r464 : std_logic_vector(0 to 0) := (others => '0');
    variable r463 : std_logic_vector(0 to 0) := (others => '0');
    variable r462 : std_logic_vector(0 to 0) := (others => '0');
    variable r461 : std_logic_vector(0 to 0) := (others => '0');
    variable r460 : std_logic_vector(0 to 0) := (others => '0');
    variable r459 : std_logic_vector(0 to 0) := (others => '0');
    variable r458 : std_logic_vector(0 to 0) := (others => '0');
    variable r457 : std_logic_vector(0 to 0) := (others => '0');
    variable r456 : std_logic_vector(0 to 0) := (others => '0');
    variable r455 : std_logic_vector(0 to 0) := (others => '0');
    variable r454 : std_logic_vector(0 to 0) := (others => '0');
    variable r453 : std_logic_vector(0 to 0) := (others => '0');
    variable r452 : std_logic_vector(0 to 0) := (others => '0');
    variable r451 : std_logic_vector(0 to 0) := (others => '0');
    variable r450 : std_logic_vector(0 to 0) := (others => '0');
    variable r449 : std_logic_vector(0 to 0) := (others => '0');
    variable r448 : std_logic_vector(0 to 0) := (others => '0');
    variable r447 : std_logic_vector(0 to 0) := (others => '0');
    variable r446 : std_logic_vector(0 to 0) := (others => '0');
    variable r445 : std_logic_vector(0 to 0) := (others => '0');
    variable r444 : std_logic_vector(0 to 0) := (others => '0');
    variable r443 : std_logic_vector(0 to 0) := (others => '0');
    variable r442 : std_logic_vector(0 to 0) := (others => '0');
    variable r441 : std_logic_vector(0 to 0) := (others => '0');
    variable r440 : std_logic_vector(0 to 0) := (others => '0');
    variable r439 : std_logic_vector(0 to 0) := (others => '0');
    variable r438 : std_logic_vector(0 to 0) := (others => '0');
    variable r437 : std_logic_vector(0 to 0) := (others => '0');
    variable r436 : std_logic_vector(0 to 0) := (others => '0');
    variable r435 : std_logic_vector(0 to 0) := (others => '0');
    variable r434 : std_logic_vector(0 to 0) := (others => '0');
    variable r433 : std_logic_vector(0 to 0) := (others => '0');
    variable r432 : std_logic_vector(0 to 0) := (others => '0');
    variable r431 : std_logic_vector(0 to 0) := (others => '0');
    variable r430 : std_logic_vector(0 to 0) := (others => '0');
    variable r429 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r430 := "0";
    null;
    r431 := (r430);
    r432 := "0";
    null;
    r433 := (r432);
    r434 := "0";
    null;
    r435 := (r434);
    r436 := "1";
    null;
    r437 := (r436);
    r438 := "1";
    null;
    r439 := (r438);
    r440 := "1";
    null;
    r441 := (r440);
    r442 := "1";
    null;
    r443 := (r442);
    r444 := "1";
    null;
    r445 := (r444);
    r446 := "1";
    null;
    r447 := (r446);
    r448 := "0";
    null;
    r449 := (r448);
    r450 := "0";
    null;
    r451 := (r450);
    r452 := "0";
    null;
    r453 := (r452);
    r454 := "0";
    null;
    r455 := (r454);
    r456 := "0";
    null;
    r457 := (r456);
    r458 := "1";
    null;
    r459 := (r458);
    r460 := "1";
    null;
    r461 := (r460);
    r462 := "1";
    null;
    r463 := (r462);
    r464 := "1";
    null;
    r465 := (r464);
    r466 := "0";
    null;
    r467 := (r466);
    r468 := "1";
    null;
    r469 := (r468);
    r470 := "1";
    null;
    r471 := (r470);
    r472 := "0";
    null;
    r473 := (r472);
    r474 := "0";
    null;
    r475 := (r474);
    r476 := "1";
    null;
    r477 := (r476);
    r478 := "1";
    null;
    r479 := (r478);
    r480 := "0";
    null;
    r481 := (r480);
    r482 := "1";
    null;
    r483 := (r482);
    r484 := "0";
    null;
    r485 := (r484);
    r486 := "1";
    null;
    r487 := (r486);
    r488 := "0";
    null;
    r489 := (r488);
    r490 := "1";
    null;
    r491 := (r490);
    r492 := "1";
    null;
    r493 := (r492);
    r429 := (r431 & r433 & r435 & r437 & r439 & r441 & r443 & r445 & r447 & r449 & r451 & r453 & r455 & r457 & r459 & r461 & r463 & r465 & r467 & r469 & r471 & r473 & r475 & r477 & r479 & r481 & r483 & r485 & r487 & r489 & r491 & r493);
    return r429;
  end rewire_MetaprogrammingRW.w1f83d9ab_428;
  function rewire_MetaprogrammingRW.w9b05688c_361 return std_logic_vector
  is
    variable r426 : std_logic_vector(0 to 0) := (others => '0');
    variable r425 : std_logic_vector(0 to 0) := (others => '0');
    variable r424 : std_logic_vector(0 to 0) := (others => '0');
    variable r423 : std_logic_vector(0 to 0) := (others => '0');
    variable r422 : std_logic_vector(0 to 0) := (others => '0');
    variable r421 : std_logic_vector(0 to 0) := (others => '0');
    variable r420 : std_logic_vector(0 to 0) := (others => '0');
    variable r419 : std_logic_vector(0 to 0) := (others => '0');
    variable r418 : std_logic_vector(0 to 0) := (others => '0');
    variable r417 : std_logic_vector(0 to 0) := (others => '0');
    variable r416 : std_logic_vector(0 to 0) := (others => '0');
    variable r415 : std_logic_vector(0 to 0) := (others => '0');
    variable r414 : std_logic_vector(0 to 0) := (others => '0');
    variable r413 : std_logic_vector(0 to 0) := (others => '0');
    variable r412 : std_logic_vector(0 to 0) := (others => '0');
    variable r411 : std_logic_vector(0 to 0) := (others => '0');
    variable r410 : std_logic_vector(0 to 0) := (others => '0');
    variable r409 : std_logic_vector(0 to 0) := (others => '0');
    variable r408 : std_logic_vector(0 to 0) := (others => '0');
    variable r407 : std_logic_vector(0 to 0) := (others => '0');
    variable r406 : std_logic_vector(0 to 0) := (others => '0');
    variable r405 : std_logic_vector(0 to 0) := (others => '0');
    variable r404 : std_logic_vector(0 to 0) := (others => '0');
    variable r403 : std_logic_vector(0 to 0) := (others => '0');
    variable r402 : std_logic_vector(0 to 0) := (others => '0');
    variable r401 : std_logic_vector(0 to 0) := (others => '0');
    variable r400 : std_logic_vector(0 to 0) := (others => '0');
    variable r399 : std_logic_vector(0 to 0) := (others => '0');
    variable r398 : std_logic_vector(0 to 0) := (others => '0');
    variable r397 : std_logic_vector(0 to 0) := (others => '0');
    variable r396 : std_logic_vector(0 to 0) := (others => '0');
    variable r395 : std_logic_vector(0 to 0) := (others => '0');
    variable r394 : std_logic_vector(0 to 0) := (others => '0');
    variable r393 : std_logic_vector(0 to 0) := (others => '0');
    variable r392 : std_logic_vector(0 to 0) := (others => '0');
    variable r391 : std_logic_vector(0 to 0) := (others => '0');
    variable r390 : std_logic_vector(0 to 0) := (others => '0');
    variable r389 : std_logic_vector(0 to 0) := (others => '0');
    variable r388 : std_logic_vector(0 to 0) := (others => '0');
    variable r387 : std_logic_vector(0 to 0) := (others => '0');
    variable r386 : std_logic_vector(0 to 0) := (others => '0');
    variable r385 : std_logic_vector(0 to 0) := (others => '0');
    variable r384 : std_logic_vector(0 to 0) := (others => '0');
    variable r383 : std_logic_vector(0 to 0) := (others => '0');
    variable r382 : std_logic_vector(0 to 0) := (others => '0');
    variable r381 : std_logic_vector(0 to 0) := (others => '0');
    variable r380 : std_logic_vector(0 to 0) := (others => '0');
    variable r379 : std_logic_vector(0 to 0) := (others => '0');
    variable r378 : std_logic_vector(0 to 0) := (others => '0');
    variable r377 : std_logic_vector(0 to 0) := (others => '0');
    variable r376 : std_logic_vector(0 to 0) := (others => '0');
    variable r375 : std_logic_vector(0 to 0) := (others => '0');
    variable r374 : std_logic_vector(0 to 0) := (others => '0');
    variable r373 : std_logic_vector(0 to 0) := (others => '0');
    variable r372 : std_logic_vector(0 to 0) := (others => '0');
    variable r371 : std_logic_vector(0 to 0) := (others => '0');
    variable r370 : std_logic_vector(0 to 0) := (others => '0');
    variable r369 : std_logic_vector(0 to 0) := (others => '0');
    variable r368 : std_logic_vector(0 to 0) := (others => '0');
    variable r367 : std_logic_vector(0 to 0) := (others => '0');
    variable r366 : std_logic_vector(0 to 0) := (others => '0');
    variable r365 : std_logic_vector(0 to 0) := (others => '0');
    variable r364 : std_logic_vector(0 to 0) := (others => '0');
    variable r363 : std_logic_vector(0 to 0) := (others => '0');
    variable r362 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r363 := "1";
    null;
    r364 := (r363);
    r365 := "0";
    null;
    r366 := (r365);
    r367 := "0";
    null;
    r368 := (r367);
    r369 := "1";
    null;
    r370 := (r369);
    r371 := "1";
    null;
    r372 := (r371);
    r373 := "0";
    null;
    r374 := (r373);
    r375 := "1";
    null;
    r376 := (r375);
    r377 := "1";
    null;
    r378 := (r377);
    r379 := "0";
    null;
    r380 := (r379);
    r381 := "0";
    null;
    r382 := (r381);
    r383 := "0";
    null;
    r384 := (r383);
    r385 := "0";
    null;
    r386 := (r385);
    r387 := "0";
    null;
    r388 := (r387);
    r389 := "1";
    null;
    r390 := (r389);
    r391 := "0";
    null;
    r392 := (r391);
    r393 := "1";
    null;
    r394 := (r393);
    r395 := "0";
    null;
    r396 := (r395);
    r397 := "1";
    null;
    r398 := (r397);
    r399 := "1";
    null;
    r400 := (r399);
    r401 := "0";
    null;
    r402 := (r401);
    r403 := "1";
    null;
    r404 := (r403);
    r405 := "0";
    null;
    r406 := (r405);
    r407 := "0";
    null;
    r408 := (r407);
    r409 := "0";
    null;
    r410 := (r409);
    r411 := "1";
    null;
    r412 := (r411);
    r413 := "0";
    null;
    r414 := (r413);
    r415 := "0";
    null;
    r416 := (r415);
    r417 := "0";
    null;
    r418 := (r417);
    r419 := "1";
    null;
    r420 := (r419);
    r421 := "1";
    null;
    r422 := (r421);
    r423 := "0";
    null;
    r424 := (r423);
    r425 := "0";
    null;
    r426 := (r425);
    r362 := (r364 & r366 & r368 & r370 & r372 & r374 & r376 & r378 & r380 & r382 & r384 & r386 & r388 & r390 & r392 & r394 & r396 & r398 & r400 & r402 & r404 & r406 & r408 & r410 & r412 & r414 & r416 & r418 & r420 & r422 & r424 & r426);
    return r362;
  end rewire_MetaprogrammingRW.w9b05688c_361;
  function rewire_MetaprogrammingRW.w510e527f_294 return std_logic_vector
  is
    variable r359 : std_logic_vector(0 to 0) := (others => '0');
    variable r358 : std_logic_vector(0 to 0) := (others => '0');
    variable r357 : std_logic_vector(0 to 0) := (others => '0');
    variable r356 : std_logic_vector(0 to 0) := (others => '0');
    variable r355 : std_logic_vector(0 to 0) := (others => '0');
    variable r354 : std_logic_vector(0 to 0) := (others => '0');
    variable r353 : std_logic_vector(0 to 0) := (others => '0');
    variable r352 : std_logic_vector(0 to 0) := (others => '0');
    variable r351 : std_logic_vector(0 to 0) := (others => '0');
    variable r350 : std_logic_vector(0 to 0) := (others => '0');
    variable r349 : std_logic_vector(0 to 0) := (others => '0');
    variable r348 : std_logic_vector(0 to 0) := (others => '0');
    variable r347 : std_logic_vector(0 to 0) := (others => '0');
    variable r346 : std_logic_vector(0 to 0) := (others => '0');
    variable r345 : std_logic_vector(0 to 0) := (others => '0');
    variable r344 : std_logic_vector(0 to 0) := (others => '0');
    variable r343 : std_logic_vector(0 to 0) := (others => '0');
    variable r342 : std_logic_vector(0 to 0) := (others => '0');
    variable r341 : std_logic_vector(0 to 0) := (others => '0');
    variable r340 : std_logic_vector(0 to 0) := (others => '0');
    variable r339 : std_logic_vector(0 to 0) := (others => '0');
    variable r338 : std_logic_vector(0 to 0) := (others => '0');
    variable r337 : std_logic_vector(0 to 0) := (others => '0');
    variable r336 : std_logic_vector(0 to 0) := (others => '0');
    variable r335 : std_logic_vector(0 to 0) := (others => '0');
    variable r334 : std_logic_vector(0 to 0) := (others => '0');
    variable r333 : std_logic_vector(0 to 0) := (others => '0');
    variable r332 : std_logic_vector(0 to 0) := (others => '0');
    variable r331 : std_logic_vector(0 to 0) := (others => '0');
    variable r330 : std_logic_vector(0 to 0) := (others => '0');
    variable r329 : std_logic_vector(0 to 0) := (others => '0');
    variable r328 : std_logic_vector(0 to 0) := (others => '0');
    variable r327 : std_logic_vector(0 to 0) := (others => '0');
    variable r326 : std_logic_vector(0 to 0) := (others => '0');
    variable r325 : std_logic_vector(0 to 0) := (others => '0');
    variable r324 : std_logic_vector(0 to 0) := (others => '0');
    variable r323 : std_logic_vector(0 to 0) := (others => '0');
    variable r322 : std_logic_vector(0 to 0) := (others => '0');
    variable r321 : std_logic_vector(0 to 0) := (others => '0');
    variable r320 : std_logic_vector(0 to 0) := (others => '0');
    variable r319 : std_logic_vector(0 to 0) := (others => '0');
    variable r318 : std_logic_vector(0 to 0) := (others => '0');
    variable r317 : std_logic_vector(0 to 0) := (others => '0');
    variable r316 : std_logic_vector(0 to 0) := (others => '0');
    variable r315 : std_logic_vector(0 to 0) := (others => '0');
    variable r314 : std_logic_vector(0 to 0) := (others => '0');
    variable r313 : std_logic_vector(0 to 0) := (others => '0');
    variable r312 : std_logic_vector(0 to 0) := (others => '0');
    variable r311 : std_logic_vector(0 to 0) := (others => '0');
    variable r310 : std_logic_vector(0 to 0) := (others => '0');
    variable r309 : std_logic_vector(0 to 0) := (others => '0');
    variable r308 : std_logic_vector(0 to 0) := (others => '0');
    variable r307 : std_logic_vector(0 to 0) := (others => '0');
    variable r306 : std_logic_vector(0 to 0) := (others => '0');
    variable r305 : std_logic_vector(0 to 0) := (others => '0');
    variable r304 : std_logic_vector(0 to 0) := (others => '0');
    variable r303 : std_logic_vector(0 to 0) := (others => '0');
    variable r302 : std_logic_vector(0 to 0) := (others => '0');
    variable r301 : std_logic_vector(0 to 0) := (others => '0');
    variable r300 : std_logic_vector(0 to 0) := (others => '0');
    variable r299 : std_logic_vector(0 to 0) := (others => '0');
    variable r298 : std_logic_vector(0 to 0) := (others => '0');
    variable r297 : std_logic_vector(0 to 0) := (others => '0');
    variable r296 : std_logic_vector(0 to 0) := (others => '0');
    variable r295 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r296 := "0";
    null;
    r297 := (r296);
    r298 := "1";
    null;
    r299 := (r298);
    r300 := "0";
    null;
    r301 := (r300);
    r302 := "1";
    null;
    r303 := (r302);
    r304 := "0";
    null;
    r305 := (r304);
    r306 := "0";
    null;
    r307 := (r306);
    r308 := "0";
    null;
    r309 := (r308);
    r310 := "1";
    null;
    r311 := (r310);
    r312 := "0";
    null;
    r313 := (r312);
    r314 := "0";
    null;
    r315 := (r314);
    r316 := "0";
    null;
    r317 := (r316);
    r318 := "0";
    null;
    r319 := (r318);
    r320 := "1";
    null;
    r321 := (r320);
    r322 := "1";
    null;
    r323 := (r322);
    r324 := "1";
    null;
    r325 := (r324);
    r326 := "0";
    null;
    r327 := (r326);
    r328 := "0";
    null;
    r329 := (r328);
    r330 := "1";
    null;
    r331 := (r330);
    r332 := "0";
    null;
    r333 := (r332);
    r334 := "1";
    null;
    r335 := (r334);
    r336 := "0";
    null;
    r337 := (r336);
    r338 := "0";
    null;
    r339 := (r338);
    r340 := "1";
    null;
    r341 := (r340);
    r342 := "0";
    null;
    r343 := (r342);
    r344 := "0";
    null;
    r345 := (r344);
    r346 := "1";
    null;
    r347 := (r346);
    r348 := "1";
    null;
    r349 := (r348);
    r350 := "1";
    null;
    r351 := (r350);
    r352 := "1";
    null;
    r353 := (r352);
    r354 := "1";
    null;
    r355 := (r354);
    r356 := "1";
    null;
    r357 := (r356);
    r358 := "1";
    null;
    r359 := (r358);
    r295 := (r297 & r299 & r301 & r303 & r305 & r307 & r309 & r311 & r313 & r315 & r317 & r319 & r321 & r323 & r325 & r327 & r329 & r331 & r333 & r335 & r337 & r339 & r341 & r343 & r345 & r347 & r349 & r351 & r353 & r355 & r357 & r359);
    return r295;
  end rewire_MetaprogrammingRW.w510e527f_294;
  function rewire_MetaprogrammingRW.wa54ff53a_227 return std_logic_vector
  is
    variable r292 : std_logic_vector(0 to 0) := (others => '0');
    variable r291 : std_logic_vector(0 to 0) := (others => '0');
    variable r290 : std_logic_vector(0 to 0) := (others => '0');
    variable r289 : std_logic_vector(0 to 0) := (others => '0');
    variable r288 : std_logic_vector(0 to 0) := (others => '0');
    variable r287 : std_logic_vector(0 to 0) := (others => '0');
    variable r286 : std_logic_vector(0 to 0) := (others => '0');
    variable r285 : std_logic_vector(0 to 0) := (others => '0');
    variable r284 : std_logic_vector(0 to 0) := (others => '0');
    variable r283 : std_logic_vector(0 to 0) := (others => '0');
    variable r282 : std_logic_vector(0 to 0) := (others => '0');
    variable r281 : std_logic_vector(0 to 0) := (others => '0');
    variable r280 : std_logic_vector(0 to 0) := (others => '0');
    variable r279 : std_logic_vector(0 to 0) := (others => '0');
    variable r278 : std_logic_vector(0 to 0) := (others => '0');
    variable r277 : std_logic_vector(0 to 0) := (others => '0');
    variable r276 : std_logic_vector(0 to 0) := (others => '0');
    variable r275 : std_logic_vector(0 to 0) := (others => '0');
    variable r274 : std_logic_vector(0 to 0) := (others => '0');
    variable r273 : std_logic_vector(0 to 0) := (others => '0');
    variable r272 : std_logic_vector(0 to 0) := (others => '0');
    variable r271 : std_logic_vector(0 to 0) := (others => '0');
    variable r270 : std_logic_vector(0 to 0) := (others => '0');
    variable r269 : std_logic_vector(0 to 0) := (others => '0');
    variable r268 : std_logic_vector(0 to 0) := (others => '0');
    variable r267 : std_logic_vector(0 to 0) := (others => '0');
    variable r266 : std_logic_vector(0 to 0) := (others => '0');
    variable r265 : std_logic_vector(0 to 0) := (others => '0');
    variable r264 : std_logic_vector(0 to 0) := (others => '0');
    variable r263 : std_logic_vector(0 to 0) := (others => '0');
    variable r262 : std_logic_vector(0 to 0) := (others => '0');
    variable r261 : std_logic_vector(0 to 0) := (others => '0');
    variable r260 : std_logic_vector(0 to 0) := (others => '0');
    variable r259 : std_logic_vector(0 to 0) := (others => '0');
    variable r258 : std_logic_vector(0 to 0) := (others => '0');
    variable r257 : std_logic_vector(0 to 0) := (others => '0');
    variable r256 : std_logic_vector(0 to 0) := (others => '0');
    variable r255 : std_logic_vector(0 to 0) := (others => '0');
    variable r254 : std_logic_vector(0 to 0) := (others => '0');
    variable r253 : std_logic_vector(0 to 0) := (others => '0');
    variable r252 : std_logic_vector(0 to 0) := (others => '0');
    variable r251 : std_logic_vector(0 to 0) := (others => '0');
    variable r250 : std_logic_vector(0 to 0) := (others => '0');
    variable r249 : std_logic_vector(0 to 0) := (others => '0');
    variable r248 : std_logic_vector(0 to 0) := (others => '0');
    variable r247 : std_logic_vector(0 to 0) := (others => '0');
    variable r246 : std_logic_vector(0 to 0) := (others => '0');
    variable r245 : std_logic_vector(0 to 0) := (others => '0');
    variable r244 : std_logic_vector(0 to 0) := (others => '0');
    variable r243 : std_logic_vector(0 to 0) := (others => '0');
    variable r242 : std_logic_vector(0 to 0) := (others => '0');
    variable r241 : std_logic_vector(0 to 0) := (others => '0');
    variable r240 : std_logic_vector(0 to 0) := (others => '0');
    variable r239 : std_logic_vector(0 to 0) := (others => '0');
    variable r238 : std_logic_vector(0 to 0) := (others => '0');
    variable r237 : std_logic_vector(0 to 0) := (others => '0');
    variable r236 : std_logic_vector(0 to 0) := (others => '0');
    variable r235 : std_logic_vector(0 to 0) := (others => '0');
    variable r234 : std_logic_vector(0 to 0) := (others => '0');
    variable r233 : std_logic_vector(0 to 0) := (others => '0');
    variable r232 : std_logic_vector(0 to 0) := (others => '0');
    variable r231 : std_logic_vector(0 to 0) := (others => '0');
    variable r230 : std_logic_vector(0 to 0) := (others => '0');
    variable r229 : std_logic_vector(0 to 0) := (others => '0');
    variable r228 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r229 := "1";
    null;
    r230 := (r229);
    r231 := "0";
    null;
    r232 := (r231);
    r233 := "1";
    null;
    r234 := (r233);
    r235 := "0";
    null;
    r236 := (r235);
    r237 := "0";
    null;
    r238 := (r237);
    r239 := "1";
    null;
    r240 := (r239);
    r241 := "0";
    null;
    r242 := (r241);
    r243 := "1";
    null;
    r244 := (r243);
    r245 := "0";
    null;
    r246 := (r245);
    r247 := "1";
    null;
    r248 := (r247);
    r249 := "0";
    null;
    r250 := (r249);
    r251 := "0";
    null;
    r252 := (r251);
    r253 := "1";
    null;
    r254 := (r253);
    r255 := "1";
    null;
    r256 := (r255);
    r257 := "1";
    null;
    r258 := (r257);
    r259 := "1";
    null;
    r260 := (r259);
    r261 := "1";
    null;
    r262 := (r261);
    r263 := "1";
    null;
    r264 := (r263);
    r265 := "1";
    null;
    r266 := (r265);
    r267 := "1";
    null;
    r268 := (r267);
    r269 := "0";
    null;
    r270 := (r269);
    r271 := "1";
    null;
    r272 := (r271);
    r273 := "0";
    null;
    r274 := (r273);
    r275 := "1";
    null;
    r276 := (r275);
    r277 := "0";
    null;
    r278 := (r277);
    r279 := "0";
    null;
    r280 := (r279);
    r281 := "1";
    null;
    r282 := (r281);
    r283 := "1";
    null;
    r284 := (r283);
    r285 := "1";
    null;
    r286 := (r285);
    r287 := "0";
    null;
    r288 := (r287);
    r289 := "1";
    null;
    r290 := (r289);
    r291 := "0";
    null;
    r292 := (r291);
    r228 := (r230 & r232 & r234 & r236 & r238 & r240 & r242 & r244 & r246 & r248 & r250 & r252 & r254 & r256 & r258 & r260 & r262 & r264 & r266 & r268 & r270 & r272 & r274 & r276 & r278 & r280 & r282 & r284 & r286 & r288 & r290 & r292);
    return r228;
  end rewire_MetaprogrammingRW.wa54ff53a_227;
  function rewire_MetaprogrammingRW.w3c6ef372_160 return std_logic_vector
  is
    variable r225 : std_logic_vector(0 to 0) := (others => '0');
    variable r224 : std_logic_vector(0 to 0) := (others => '0');
    variable r223 : std_logic_vector(0 to 0) := (others => '0');
    variable r222 : std_logic_vector(0 to 0) := (others => '0');
    variable r221 : std_logic_vector(0 to 0) := (others => '0');
    variable r220 : std_logic_vector(0 to 0) := (others => '0');
    variable r219 : std_logic_vector(0 to 0) := (others => '0');
    variable r218 : std_logic_vector(0 to 0) := (others => '0');
    variable r217 : std_logic_vector(0 to 0) := (others => '0');
    variable r216 : std_logic_vector(0 to 0) := (others => '0');
    variable r215 : std_logic_vector(0 to 0) := (others => '0');
    variable r214 : std_logic_vector(0 to 0) := (others => '0');
    variable r213 : std_logic_vector(0 to 0) := (others => '0');
    variable r212 : std_logic_vector(0 to 0) := (others => '0');
    variable r211 : std_logic_vector(0 to 0) := (others => '0');
    variable r210 : std_logic_vector(0 to 0) := (others => '0');
    variable r209 : std_logic_vector(0 to 0) := (others => '0');
    variable r208 : std_logic_vector(0 to 0) := (others => '0');
    variable r207 : std_logic_vector(0 to 0) := (others => '0');
    variable r206 : std_logic_vector(0 to 0) := (others => '0');
    variable r205 : std_logic_vector(0 to 0) := (others => '0');
    variable r204 : std_logic_vector(0 to 0) := (others => '0');
    variable r203 : std_logic_vector(0 to 0) := (others => '0');
    variable r202 : std_logic_vector(0 to 0) := (others => '0');
    variable r201 : std_logic_vector(0 to 0) := (others => '0');
    variable r200 : std_logic_vector(0 to 0) := (others => '0');
    variable r199 : std_logic_vector(0 to 0) := (others => '0');
    variable r198 : std_logic_vector(0 to 0) := (others => '0');
    variable r197 : std_logic_vector(0 to 0) := (others => '0');
    variable r196 : std_logic_vector(0 to 0) := (others => '0');
    variable r195 : std_logic_vector(0 to 0) := (others => '0');
    variable r194 : std_logic_vector(0 to 0) := (others => '0');
    variable r193 : std_logic_vector(0 to 0) := (others => '0');
    variable r192 : std_logic_vector(0 to 0) := (others => '0');
    variable r191 : std_logic_vector(0 to 0) := (others => '0');
    variable r190 : std_logic_vector(0 to 0) := (others => '0');
    variable r189 : std_logic_vector(0 to 0) := (others => '0');
    variable r188 : std_logic_vector(0 to 0) := (others => '0');
    variable r187 : std_logic_vector(0 to 0) := (others => '0');
    variable r186 : std_logic_vector(0 to 0) := (others => '0');
    variable r185 : std_logic_vector(0 to 0) := (others => '0');
    variable r184 : std_logic_vector(0 to 0) := (others => '0');
    variable r183 : std_logic_vector(0 to 0) := (others => '0');
    variable r182 : std_logic_vector(0 to 0) := (others => '0');
    variable r181 : std_logic_vector(0 to 0) := (others => '0');
    variable r180 : std_logic_vector(0 to 0) := (others => '0');
    variable r179 : std_logic_vector(0 to 0) := (others => '0');
    variable r178 : std_logic_vector(0 to 0) := (others => '0');
    variable r177 : std_logic_vector(0 to 0) := (others => '0');
    variable r176 : std_logic_vector(0 to 0) := (others => '0');
    variable r175 : std_logic_vector(0 to 0) := (others => '0');
    variable r174 : std_logic_vector(0 to 0) := (others => '0');
    variable r173 : std_logic_vector(0 to 0) := (others => '0');
    variable r172 : std_logic_vector(0 to 0) := (others => '0');
    variable r171 : std_logic_vector(0 to 0) := (others => '0');
    variable r170 : std_logic_vector(0 to 0) := (others => '0');
    variable r169 : std_logic_vector(0 to 0) := (others => '0');
    variable r168 : std_logic_vector(0 to 0) := (others => '0');
    variable r167 : std_logic_vector(0 to 0) := (others => '0');
    variable r166 : std_logic_vector(0 to 0) := (others => '0');
    variable r165 : std_logic_vector(0 to 0) := (others => '0');
    variable r164 : std_logic_vector(0 to 0) := (others => '0');
    variable r163 : std_logic_vector(0 to 0) := (others => '0');
    variable r162 : std_logic_vector(0 to 0) := (others => '0');
    variable r161 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r162 := "0";
    null;
    r163 := (r162);
    r164 := "0";
    null;
    r165 := (r164);
    r166 := "1";
    null;
    r167 := (r166);
    r168 := "1";
    null;
    r169 := (r168);
    r170 := "1";
    null;
    r171 := (r170);
    r172 := "1";
    null;
    r173 := (r172);
    r174 := "0";
    null;
    r175 := (r174);
    r176 := "0";
    null;
    r177 := (r176);
    r178 := "0";
    null;
    r179 := (r178);
    r180 := "1";
    null;
    r181 := (r180);
    r182 := "1";
    null;
    r183 := (r182);
    r184 := "0";
    null;
    r185 := (r184);
    r186 := "1";
    null;
    r187 := (r186);
    r188 := "1";
    null;
    r189 := (r188);
    r190 := "1";
    null;
    r191 := (r190);
    r192 := "0";
    null;
    r193 := (r192);
    r194 := "1";
    null;
    r195 := (r194);
    r196 := "1";
    null;
    r197 := (r196);
    r198 := "1";
    null;
    r199 := (r198);
    r200 := "1";
    null;
    r201 := (r200);
    r202 := "0";
    null;
    r203 := (r202);
    r204 := "0";
    null;
    r205 := (r204);
    r206 := "1";
    null;
    r207 := (r206);
    r208 := "1";
    null;
    r209 := (r208);
    r210 := "0";
    null;
    r211 := (r210);
    r212 := "1";
    null;
    r213 := (r212);
    r214 := "1";
    null;
    r215 := (r214);
    r216 := "1";
    null;
    r217 := (r216);
    r218 := "0";
    null;
    r219 := (r218);
    r220 := "0";
    null;
    r221 := (r220);
    r222 := "1";
    null;
    r223 := (r222);
    r224 := "0";
    null;
    r225 := (r224);
    r161 := (r163 & r165 & r167 & r169 & r171 & r173 & r175 & r177 & r179 & r181 & r183 & r185 & r187 & r189 & r191 & r193 & r195 & r197 & r199 & r201 & r203 & r205 & r207 & r209 & r211 & r213 & r215 & r217 & r219 & r221 & r223 & r225);
    return r161;
  end rewire_MetaprogrammingRW.w3c6ef372_160;
  function rewire_MetaprogrammingRW.wbb67ae85_93 return std_logic_vector
  is
    variable r158 : std_logic_vector(0 to 0) := (others => '0');
    variable r157 : std_logic_vector(0 to 0) := (others => '0');
    variable r156 : std_logic_vector(0 to 0) := (others => '0');
    variable r155 : std_logic_vector(0 to 0) := (others => '0');
    variable r154 : std_logic_vector(0 to 0) := (others => '0');
    variable r153 : std_logic_vector(0 to 0) := (others => '0');
    variable r152 : std_logic_vector(0 to 0) := (others => '0');
    variable r151 : std_logic_vector(0 to 0) := (others => '0');
    variable r150 : std_logic_vector(0 to 0) := (others => '0');
    variable r149 : std_logic_vector(0 to 0) := (others => '0');
    variable r148 : std_logic_vector(0 to 0) := (others => '0');
    variable r147 : std_logic_vector(0 to 0) := (others => '0');
    variable r146 : std_logic_vector(0 to 0) := (others => '0');
    variable r145 : std_logic_vector(0 to 0) := (others => '0');
    variable r144 : std_logic_vector(0 to 0) := (others => '0');
    variable r143 : std_logic_vector(0 to 0) := (others => '0');
    variable r142 : std_logic_vector(0 to 0) := (others => '0');
    variable r141 : std_logic_vector(0 to 0) := (others => '0');
    variable r140 : std_logic_vector(0 to 0) := (others => '0');
    variable r139 : std_logic_vector(0 to 0) := (others => '0');
    variable r138 : std_logic_vector(0 to 0) := (others => '0');
    variable r137 : std_logic_vector(0 to 0) := (others => '0');
    variable r136 : std_logic_vector(0 to 0) := (others => '0');
    variable r135 : std_logic_vector(0 to 0) := (others => '0');
    variable r134 : std_logic_vector(0 to 0) := (others => '0');
    variable r133 : std_logic_vector(0 to 0) := (others => '0');
    variable r132 : std_logic_vector(0 to 0) := (others => '0');
    variable r131 : std_logic_vector(0 to 0) := (others => '0');
    variable r130 : std_logic_vector(0 to 0) := (others => '0');
    variable r129 : std_logic_vector(0 to 0) := (others => '0');
    variable r128 : std_logic_vector(0 to 0) := (others => '0');
    variable r127 : std_logic_vector(0 to 0) := (others => '0');
    variable r126 : std_logic_vector(0 to 0) := (others => '0');
    variable r125 : std_logic_vector(0 to 0) := (others => '0');
    variable r124 : std_logic_vector(0 to 0) := (others => '0');
    variable r123 : std_logic_vector(0 to 0) := (others => '0');
    variable r122 : std_logic_vector(0 to 0) := (others => '0');
    variable r121 : std_logic_vector(0 to 0) := (others => '0');
    variable r120 : std_logic_vector(0 to 0) := (others => '0');
    variable r119 : std_logic_vector(0 to 0) := (others => '0');
    variable r118 : std_logic_vector(0 to 0) := (others => '0');
    variable r117 : std_logic_vector(0 to 0) := (others => '0');
    variable r116 : std_logic_vector(0 to 0) := (others => '0');
    variable r115 : std_logic_vector(0 to 0) := (others => '0');
    variable r114 : std_logic_vector(0 to 0) := (others => '0');
    variable r113 : std_logic_vector(0 to 0) := (others => '0');
    variable r112 : std_logic_vector(0 to 0) := (others => '0');
    variable r111 : std_logic_vector(0 to 0) := (others => '0');
    variable r110 : std_logic_vector(0 to 0) := (others => '0');
    variable r109 : std_logic_vector(0 to 0) := (others => '0');
    variable r108 : std_logic_vector(0 to 0) := (others => '0');
    variable r107 : std_logic_vector(0 to 0) := (others => '0');
    variable r106 : std_logic_vector(0 to 0) := (others => '0');
    variable r105 : std_logic_vector(0 to 0) := (others => '0');
    variable r104 : std_logic_vector(0 to 0) := (others => '0');
    variable r103 : std_logic_vector(0 to 0) := (others => '0');
    variable r102 : std_logic_vector(0 to 0) := (others => '0');
    variable r101 : std_logic_vector(0 to 0) := (others => '0');
    variable r100 : std_logic_vector(0 to 0) := (others => '0');
    variable r99 : std_logic_vector(0 to 0) := (others => '0');
    variable r98 : std_logic_vector(0 to 0) := (others => '0');
    variable r97 : std_logic_vector(0 to 0) := (others => '0');
    variable r96 : std_logic_vector(0 to 0) := (others => '0');
    variable r95 : std_logic_vector(0 to 0) := (others => '0');
    variable r94 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r95 := "1";
    null;
    r96 := (r95);
    r97 := "0";
    null;
    r98 := (r97);
    r99 := "1";
    null;
    r100 := (r99);
    r101 := "1";
    null;
    r102 := (r101);
    r103 := "1";
    null;
    r104 := (r103);
    r105 := "0";
    null;
    r106 := (r105);
    r107 := "1";
    null;
    r108 := (r107);
    r109 := "1";
    null;
    r110 := (r109);
    r111 := "0";
    null;
    r112 := (r111);
    r113 := "1";
    null;
    r114 := (r113);
    r115 := "1";
    null;
    r116 := (r115);
    r117 := "0";
    null;
    r118 := (r117);
    r119 := "0";
    null;
    r120 := (r119);
    r121 := "1";
    null;
    r122 := (r121);
    r123 := "1";
    null;
    r124 := (r123);
    r125 := "1";
    null;
    r126 := (r125);
    r127 := "1";
    null;
    r128 := (r127);
    r129 := "0";
    null;
    r130 := (r129);
    r131 := "1";
    null;
    r132 := (r131);
    r133 := "0";
    null;
    r134 := (r133);
    r135 := "1";
    null;
    r136 := (r135);
    r137 := "1";
    null;
    r138 := (r137);
    r139 := "1";
    null;
    r140 := (r139);
    r141 := "0";
    null;
    r142 := (r141);
    r143 := "1";
    null;
    r144 := (r143);
    r145 := "0";
    null;
    r146 := (r145);
    r147 := "0";
    null;
    r148 := (r147);
    r149 := "0";
    null;
    r150 := (r149);
    r151 := "0";
    null;
    r152 := (r151);
    r153 := "1";
    null;
    r154 := (r153);
    r155 := "0";
    null;
    r156 := (r155);
    r157 := "1";
    null;
    r158 := (r157);
    r94 := (r96 & r98 & r100 & r102 & r104 & r106 & r108 & r110 & r112 & r114 & r116 & r118 & r120 & r122 & r124 & r126 & r128 & r130 & r132 & r134 & r136 & r138 & r140 & r142 & r144 & r146 & r148 & r150 & r152 & r154 & r156 & r158);
    return r94;
  end rewire_MetaprogrammingRW.wbb67ae85_93;
  function rewire_MetaprogrammingRW.w6a09e667_26 return std_logic_vector
  is
    variable r91 : std_logic_vector(0 to 0) := (others => '0');
    variable r90 : std_logic_vector(0 to 0) := (others => '0');
    variable r89 : std_logic_vector(0 to 0) := (others => '0');
    variable r88 : std_logic_vector(0 to 0) := (others => '0');
    variable r87 : std_logic_vector(0 to 0) := (others => '0');
    variable r86 : std_logic_vector(0 to 0) := (others => '0');
    variable r85 : std_logic_vector(0 to 0) := (others => '0');
    variable r84 : std_logic_vector(0 to 0) := (others => '0');
    variable r83 : std_logic_vector(0 to 0) := (others => '0');
    variable r82 : std_logic_vector(0 to 0) := (others => '0');
    variable r81 : std_logic_vector(0 to 0) := (others => '0');
    variable r80 : std_logic_vector(0 to 0) := (others => '0');
    variable r79 : std_logic_vector(0 to 0) := (others => '0');
    variable r78 : std_logic_vector(0 to 0) := (others => '0');
    variable r77 : std_logic_vector(0 to 0) := (others => '0');
    variable r76 : std_logic_vector(0 to 0) := (others => '0');
    variable r75 : std_logic_vector(0 to 0) := (others => '0');
    variable r74 : std_logic_vector(0 to 0) := (others => '0');
    variable r73 : std_logic_vector(0 to 0) := (others => '0');
    variable r72 : std_logic_vector(0 to 0) := (others => '0');
    variable r71 : std_logic_vector(0 to 0) := (others => '0');
    variable r70 : std_logic_vector(0 to 0) := (others => '0');
    variable r69 : std_logic_vector(0 to 0) := (others => '0');
    variable r68 : std_logic_vector(0 to 0) := (others => '0');
    variable r67 : std_logic_vector(0 to 0) := (others => '0');
    variable r66 : std_logic_vector(0 to 0) := (others => '0');
    variable r65 : std_logic_vector(0 to 0) := (others => '0');
    variable r64 : std_logic_vector(0 to 0) := (others => '0');
    variable r63 : std_logic_vector(0 to 0) := (others => '0');
    variable r62 : std_logic_vector(0 to 0) := (others => '0');
    variable r61 : std_logic_vector(0 to 0) := (others => '0');
    variable r60 : std_logic_vector(0 to 0) := (others => '0');
    variable r59 : std_logic_vector(0 to 0) := (others => '0');
    variable r58 : std_logic_vector(0 to 0) := (others => '0');
    variable r57 : std_logic_vector(0 to 0) := (others => '0');
    variable r56 : std_logic_vector(0 to 0) := (others => '0');
    variable r55 : std_logic_vector(0 to 0) := (others => '0');
    variable r54 : std_logic_vector(0 to 0) := (others => '0');
    variable r53 : std_logic_vector(0 to 0) := (others => '0');
    variable r52 : std_logic_vector(0 to 0) := (others => '0');
    variable r51 : std_logic_vector(0 to 0) := (others => '0');
    variable r50 : std_logic_vector(0 to 0) := (others => '0');
    variable r49 : std_logic_vector(0 to 0) := (others => '0');
    variable r48 : std_logic_vector(0 to 0) := (others => '0');
    variable r47 : std_logic_vector(0 to 0) := (others => '0');
    variable r46 : std_logic_vector(0 to 0) := (others => '0');
    variable r45 : std_logic_vector(0 to 0) := (others => '0');
    variable r44 : std_logic_vector(0 to 0) := (others => '0');
    variable r43 : std_logic_vector(0 to 0) := (others => '0');
    variable r42 : std_logic_vector(0 to 0) := (others => '0');
    variable r41 : std_logic_vector(0 to 0) := (others => '0');
    variable r40 : std_logic_vector(0 to 0) := (others => '0');
    variable r39 : std_logic_vector(0 to 0) := (others => '0');
    variable r38 : std_logic_vector(0 to 0) := (others => '0');
    variable r37 : std_logic_vector(0 to 0) := (others => '0');
    variable r36 : std_logic_vector(0 to 0) := (others => '0');
    variable r35 : std_logic_vector(0 to 0) := (others => '0');
    variable r34 : std_logic_vector(0 to 0) := (others => '0');
    variable r33 : std_logic_vector(0 to 0) := (others => '0');
    variable r32 : std_logic_vector(0 to 0) := (others => '0');
    variable r31 : std_logic_vector(0 to 0) := (others => '0');
    variable r30 : std_logic_vector(0 to 0) := (others => '0');
    variable r29 : std_logic_vector(0 to 0) := (others => '0');
    variable r28 : std_logic_vector(0 to 0) := (others => '0');
    variable r27 : std_logic_vector(0 to 31) := (others => '0');
  begin
    null;
    null;
    r28 := "0";
    null;
    r29 := (r28);
    r30 := "1";
    null;
    r31 := (r30);
    r32 := "1";
    null;
    r33 := (r32);
    r34 := "0";
    null;
    r35 := (r34);
    r36 := "1";
    null;
    r37 := (r36);
    r38 := "0";
    null;
    r39 := (r38);
    r40 := "1";
    null;
    r41 := (r40);
    r42 := "0";
    null;
    r43 := (r42);
    r44 := "0";
    null;
    r45 := (r44);
    r46 := "0";
    null;
    r47 := (r46);
    r48 := "0";
    null;
    r49 := (r48);
    r50 := "0";
    null;
    r51 := (r50);
    r52 := "1";
    null;
    r53 := (r52);
    r54 := "0";
    null;
    r55 := (r54);
    r56 := "0";
    null;
    r57 := (r56);
    r58 := "1";
    null;
    r59 := (r58);
    r60 := "1";
    null;
    r61 := (r60);
    r62 := "1";
    null;
    r63 := (r62);
    r64 := "1";
    null;
    r65 := (r64);
    r66 := "0";
    null;
    r67 := (r66);
    r68 := "0";
    null;
    r69 := (r68);
    r70 := "1";
    null;
    r71 := (r70);
    r72 := "1";
    null;
    r73 := (r72);
    r74 := "0";
    null;
    r75 := (r74);
    r76 := "0";
    null;
    r77 := (r76);
    r78 := "1";
    null;
    r79 := (r78);
    r80 := "1";
    null;
    r81 := (r80);
    r82 := "0";
    null;
    r83 := (r82);
    r84 := "0";
    null;
    r85 := (r84);
    r86 := "1";
    null;
    r87 := (r86);
    r88 := "1";
    null;
    r89 := (r88);
    r90 := "1";
    null;
    r91 := (r90);
    r27 := (r29 & r31 & r33 & r35 & r37 & r39 & r41 & r43 & r45 & r47 & r49 & r51 & r53 & r55 & r57 & r59 & r61 & r63 & r65 & r67 & r69 & r71 & r73 & r75 & r77 & r79 & r81 & r83 & r85 & r87 & r89 & r91);
    return r27;
  end rewire_MetaprogrammingRW.w6a09e667_26;
  signal control_flop : control_state := STATE0;
  signal control_flop_next : control_state := STATE0;
  signal input_flop : std_logic_vector(0 to 513) := (others => '0');
  signal goto_L6287_flop : boolean := false;
  signal goto_L6280_flop : boolean := false;
  signal goto_L6264_flop : boolean := false;
  signal goto_L6110_flop : boolean := false;
  signal goto_L6230_flop : boolean := false;
  signal goto_L6115_flop : boolean := false;
  signal goto_L585_flop : boolean := false;
  signal goto_L586_flop : boolean := false;
  signal goto_L11_flop : boolean := false;
  signal goto_L13_flop : boolean := false;
  signal goto_L6233_flop : boolean := false;
  signal goto_L6266_flop : boolean := false;
  signal goto_L6245_flop : boolean := false;
  signal goto_L563_flop : boolean := false;
  signal goto_L0_flop : boolean := false;
  signal goto_L6288_flop : boolean := false;
  signal r6279_flop : std_logic_vector(0 to 513) := (others => '0');
  signal r6274_flop : std_logic_vector(0 to 257) := (others => '0');
  signal r6272_flop : std_logic_vector(0 to 1) := (others => '0');
  signal r6270_flop : std_logic_vector(0 to 255) := (others => '0');
  signal r6263_flop : std_logic_vector(0 to 513) := (others => '0');
  signal r6259_flop : std_logic_vector(0 to 255) := (others => '0');
  signal r6258_flop : std_logic_vector(0 to 257) := (others => '0');
  signal r6256_flop : std_logic_vector(0 to 1) := (others => '0');
  signal r6250_flop : std_logic_vector(0 to 5) := (others => '0');
  signal r6248_flop : std_logic_vector(0 to 5) := (others => '0');
  signal r6244_flop : std_logic_vector(0 to 255) := (others => '0');
  signal b6242_flop : boolean := false;
  signal b6240_flop : boolean := false;
  signal r6238_flop : std_logic_vector(0 to 511) := (others => '0');
  signal b6236_flop : boolean := false;
  signal r6219_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r6215_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r6211_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r6207_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r6203_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r6199_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r6195_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r6191_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r6187_flop : std_logic_vector(0 to 255) := (others => '0');
  signal b6184_flop : boolean := false;
  signal b6182_flop : boolean := false;
  signal b6180_flop : boolean := false;
  signal b6178_flop : boolean := false;
  signal b6176_flop : boolean := false;
  signal b6174_flop : boolean := false;
  signal b6172_flop : boolean := false;
  signal b6170_flop : boolean := false;
  signal r6168_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r6166_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r6164_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r6162_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r6160_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r6158_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r6156_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r6154_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r6150_flop : std_logic_vector(0 to 255) := (others => '0');
  signal b6148_flop : boolean := false;
  signal b6146_flop : boolean := false;
  signal b6144_flop : boolean := false;
  signal b6142_flop : boolean := false;
  signal b6140_flop : boolean := false;
  signal b6138_flop : boolean := false;
  signal b6136_flop : boolean := false;
  signal b6134_flop : boolean := false;
  signal r6132_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r6130_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r6128_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r6126_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r6124_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r6122_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r6120_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r6118_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r6114_flop : std_logic_vector(0 to 255) := (others => '0');
  signal b6112_flop : boolean := false;
  signal r6109_flop : std_logic_vector(0 to 513) := (others => '0');
  signal r6105_flop : std_logic_vector(0 to 255) := (others => '0');
  signal r6104_flop : std_logic_vector(0 to 257) := (others => '0');
  signal r6102_flop : std_logic_vector(0 to 1) := (others => '0');
  signal r6098_flop : std_logic_vector(0 to 5) := (others => '0');
  signal r6094_flop : std_logic_vector(0 to 255) := (others => '0');
  signal r6090_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1672_flop : std_logic_vector(0 to 5) := (others => '0');
  signal r1174_flop : std_logic_vector(0 to 255) := (others => '0');
  signal r1173_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1172_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r1169_flop : std_logic_vector(0 to 255) := (others => '0');
  signal r1163_flop : std_logic_vector(0 to 511) := (others => '0');
  signal r660_flop : std_logic_vector(0 to 511) := (others => '0');
  signal b657_flop : boolean := false;
  signal b655_flop : boolean := false;
  signal b653_flop : boolean := false;
  signal b651_flop : boolean := false;
  signal b649_flop : boolean := false;
  signal b647_flop : boolean := false;
  signal b645_flop : boolean := false;
  signal b643_flop : boolean := false;
  signal b641_flop : boolean := false;
  signal b639_flop : boolean := false;
  signal b637_flop : boolean := false;
  signal b635_flop : boolean := false;
  signal b633_flop : boolean := false;
  signal b631_flop : boolean := false;
  signal b629_flop : boolean := false;
  signal b627_flop : boolean := false;
  signal r625_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r623_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r621_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r619_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r617_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r615_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r613_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r611_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r609_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r607_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r605_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r603_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r601_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r599_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r597_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r595_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r593_flop : std_logic_vector(0 to 31) := (others => '0');
  signal r590_flop : std_logic_vector(0 to 511) := (others => '0');
  signal r588_flop : std_logic_vector(0 to 5) := (others => '0');
  signal r584_flop : std_logic_vector(0 to 513) := (others => '0');
  signal r580_flop : std_logic_vector(0 to 255) := (others => '0');
  signal r579_flop : std_logic_vector(0 to 257) := (others => '0');
  signal r577_flop : std_logic_vector(0 to 1) := (others => '0');
  signal r571_flop : std_logic_vector(0 to 255) := (others => '0');
  signal r567_flop : std_logic_vector(0 to 5) := (others => '0');
  signal r565_flop : std_logic_vector(0 to 5) := (others => '0');
  signal r562_flop : std_logic_vector(0 to 255) := (others => '0');
  signal b22_flop : boolean := false;
  signal b20_flop : boolean := false;
  signal r18_flop : std_logic_vector(0 to 511) := (others => '0');
  signal b16_flop : boolean := false;
  signal r12_flop : std_logic_vector(0 to 513) := (others => '0');
  signal r10_flop : std_logic_vector(0 to 513) := (others => '0');
  signal r6_flop : std_logic_vector(0 to 255) := (others => '0');
  signal r5_flop : std_logic_vector(0 to 257) := (others => '0');
  signal r3_flop : std_logic_vector(0 to 1) := (others => '0');
  signal statevar0_flop : std_logic_vector(0 to 255) := (others => '0');
  signal statevar1_flop : std_logic_vector(0 to 511) := (others => '0');
  signal statevar2_flop : std_logic_vector(0 to 255) := (others => '0');
  signal statevar3_flop : std_logic_vector(0 to 5) := (others => '0');
  signal goto_L6287_flop_next : boolean := false;
  signal goto_L6280_flop_next : boolean := false;
  signal goto_L6264_flop_next : boolean := false;
  signal goto_L6110_flop_next : boolean := false;
  signal goto_L6230_flop_next : boolean := false;
  signal goto_L6115_flop_next : boolean := false;
  signal goto_L585_flop_next : boolean := false;
  signal goto_L586_flop_next : boolean := false;
  signal goto_L11_flop_next : boolean := false;
  signal goto_L13_flop_next : boolean := false;
  signal goto_L6233_flop_next : boolean := false;
  signal goto_L6266_flop_next : boolean := false;
  signal goto_L6245_flop_next : boolean := false;
  signal goto_L563_flop_next : boolean := false;
  signal goto_L0_flop_next : boolean := false;
  signal goto_L6288_flop_next : boolean := false;
  signal r6279_flop_next : std_logic_vector(0 to 513) := (others => '0');
  signal r6274_flop_next : std_logic_vector(0 to 257) := (others => '0');
  signal r6272_flop_next : std_logic_vector(0 to 1) := (others => '0');
  signal r6270_flop_next : std_logic_vector(0 to 255) := (others => '0');
  signal r6263_flop_next : std_logic_vector(0 to 513) := (others => '0');
  signal r6259_flop_next : std_logic_vector(0 to 255) := (others => '0');
  signal r6258_flop_next : std_logic_vector(0 to 257) := (others => '0');
  signal r6256_flop_next : std_logic_vector(0 to 1) := (others => '0');
  signal r6250_flop_next : std_logic_vector(0 to 5) := (others => '0');
  signal r6248_flop_next : std_logic_vector(0 to 5) := (others => '0');
  signal r6244_flop_next : std_logic_vector(0 to 255) := (others => '0');
  signal b6242_flop_next : boolean := false;
  signal b6240_flop_next : boolean := false;
  signal r6238_flop_next : std_logic_vector(0 to 511) := (others => '0');
  signal b6236_flop_next : boolean := false;
  signal r6219_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r6215_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r6211_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r6207_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r6203_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r6199_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r6195_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r6191_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r6187_flop_next : std_logic_vector(0 to 255) := (others => '0');
  signal b6184_flop_next : boolean := false;
  signal b6182_flop_next : boolean := false;
  signal b6180_flop_next : boolean := false;
  signal b6178_flop_next : boolean := false;
  signal b6176_flop_next : boolean := false;
  signal b6174_flop_next : boolean := false;
  signal b6172_flop_next : boolean := false;
  signal b6170_flop_next : boolean := false;
  signal r6168_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r6166_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r6164_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r6162_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r6160_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r6158_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r6156_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r6154_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r6150_flop_next : std_logic_vector(0 to 255) := (others => '0');
  signal b6148_flop_next : boolean := false;
  signal b6146_flop_next : boolean := false;
  signal b6144_flop_next : boolean := false;
  signal b6142_flop_next : boolean := false;
  signal b6140_flop_next : boolean := false;
  signal b6138_flop_next : boolean := false;
  signal b6136_flop_next : boolean := false;
  signal b6134_flop_next : boolean := false;
  signal r6132_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r6130_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r6128_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r6126_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r6124_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r6122_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r6120_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r6118_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r6114_flop_next : std_logic_vector(0 to 255) := (others => '0');
  signal b6112_flop_next : boolean := false;
  signal r6109_flop_next : std_logic_vector(0 to 513) := (others => '0');
  signal r6105_flop_next : std_logic_vector(0 to 255) := (others => '0');
  signal r6104_flop_next : std_logic_vector(0 to 257) := (others => '0');
  signal r6102_flop_next : std_logic_vector(0 to 1) := (others => '0');
  signal r6098_flop_next : std_logic_vector(0 to 5) := (others => '0');
  signal r6094_flop_next : std_logic_vector(0 to 255) := (others => '0');
  signal r6090_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1672_flop_next : std_logic_vector(0 to 5) := (others => '0');
  signal r1174_flop_next : std_logic_vector(0 to 255) := (others => '0');
  signal r1173_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1172_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r1169_flop_next : std_logic_vector(0 to 255) := (others => '0');
  signal r1163_flop_next : std_logic_vector(0 to 511) := (others => '0');
  signal r660_flop_next : std_logic_vector(0 to 511) := (others => '0');
  signal b657_flop_next : boolean := false;
  signal b655_flop_next : boolean := false;
  signal b653_flop_next : boolean := false;
  signal b651_flop_next : boolean := false;
  signal b649_flop_next : boolean := false;
  signal b647_flop_next : boolean := false;
  signal b645_flop_next : boolean := false;
  signal b643_flop_next : boolean := false;
  signal b641_flop_next : boolean := false;
  signal b639_flop_next : boolean := false;
  signal b637_flop_next : boolean := false;
  signal b635_flop_next : boolean := false;
  signal b633_flop_next : boolean := false;
  signal b631_flop_next : boolean := false;
  signal b629_flop_next : boolean := false;
  signal b627_flop_next : boolean := false;
  signal r625_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r623_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r621_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r619_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r617_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r615_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r613_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r611_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r609_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r607_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r605_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r603_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r601_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r599_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r597_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r595_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r593_flop_next : std_logic_vector(0 to 31) := (others => '0');
  signal r590_flop_next : std_logic_vector(0 to 511) := (others => '0');
  signal r588_flop_next : std_logic_vector(0 to 5) := (others => '0');
  signal r584_flop_next : std_logic_vector(0 to 513) := (others => '0');
  signal r580_flop_next : std_logic_vector(0 to 255) := (others => '0');
  signal r579_flop_next : std_logic_vector(0 to 257) := (others => '0');
  signal r577_flop_next : std_logic_vector(0 to 1) := (others => '0');
  signal r571_flop_next : std_logic_vector(0 to 255) := (others => '0');
  signal r567_flop_next : std_logic_vector(0 to 5) := (others => '0');
  signal r565_flop_next : std_logic_vector(0 to 5) := (others => '0');
  signal r562_flop_next : std_logic_vector(0 to 255) := (others => '0');
  signal b22_flop_next : boolean := false;
  signal b20_flop_next : boolean := false;
  signal r18_flop_next : std_logic_vector(0 to 511) := (others => '0');
  signal b16_flop_next : boolean := false;
  signal r12_flop_next : std_logic_vector(0 to 513) := (others => '0');
  signal r10_flop_next : std_logic_vector(0 to 513) := (others => '0');
  signal r6_flop_next : std_logic_vector(0 to 255) := (others => '0');
  signal r5_flop_next : std_logic_vector(0 to 257) := (others => '0');
  signal r3_flop_next : std_logic_vector(0 to 1) := (others => '0');
  signal statevar0_flop_next : std_logic_vector(0 to 255) := (others => '0');
  signal statevar1_flop_next : std_logic_vector(0 to 511) := (others => '0');
  signal statevar2_flop_next : std_logic_vector(0 to 255) := (others => '0');
  signal statevar3_flop_next : std_logic_vector(0 to 5) := (others => '0');
begin
  -- Logic loop process.
  process (control_flop,input_flop,goto_L6287_flop,goto_L6280_flop,goto_L6264_flop,goto_L6110_flop,goto_L6230_flop,goto_L6115_flop,goto_L585_flop,goto_L586_flop,goto_L11_flop,goto_L13_flop,goto_L6233_flop,goto_L6266_flop,goto_L6245_flop,goto_L563_flop,goto_L0_flop,goto_L6288_flop,r6279_flop,r6274_flop,r6272_flop,r6270_flop,r6263_flop,r6259_flop,r6258_flop,r6256_flop,r6250_flop,r6248_flop,r6244_flop,b6242_flop,b6240_flop,r6238_flop,b6236_flop,r6219_flop,r6215_flop,r6211_flop,r6207_flop,r6203_flop,r6199_flop,r6195_flop,r6191_flop,r6187_flop,b6184_flop,b6182_flop,b6180_flop,b6178_flop,b6176_flop,b6174_flop,b6172_flop,b6170_flop,r6168_flop,r6166_flop,r6164_flop,r6162_flop,r6160_flop,r6158_flop,r6156_flop,r6154_flop,r6150_flop,b6148_flop,b6146_flop,b6144_flop,b6142_flop,b6140_flop,b6138_flop,b6136_flop,b6134_flop,r6132_flop,r6130_flop,r6128_flop,r6126_flop,r6124_flop,r6122_flop,r6120_flop,r6118_flop,r6114_flop,b6112_flop,r6109_flop,r6105_flop,r6104_flop,r6102_flop,r6098_flop,r6094_flop,r6090_flop,r1672_flop,r1174_flop,r1173_flop,r1172_flop,r1169_flop,r1163_flop,r660_flop,b657_flop,b655_flop,b653_flop,b651_flop,b649_flop,b647_flop,b645_flop,b643_flop,b641_flop,b639_flop,b637_flop,b635_flop,b633_flop,b631_flop,b629_flop,b627_flop,r625_flop,r623_flop,r621_flop,r619_flop,r617_flop,r615_flop,r613_flop,r611_flop,r609_flop,r607_flop,r605_flop,r603_flop,r601_flop,r599_flop,r597_flop,r595_flop,r593_flop,r590_flop,r588_flop,r584_flop,r580_flop,r579_flop,r577_flop,r571_flop,r567_flop,r565_flop,r562_flop,b22_flop,b20_flop,r18_flop,b16_flop,r12_flop,r10_flop,r6_flop,r5_flop,r3_flop,statevar0_flop,statevar1_flop,statevar2_flop,statevar3_flop)
    variable control : control_state;
    variable input_tmp : std_logic_vector(0 to 513);
    variable goto_L6287 : boolean := false;
    variable goto_L6280 : boolean := false;
    variable goto_L6264 : boolean := false;
    variable goto_L6110 : boolean := false;
    variable goto_L6230 : boolean := false;
    variable goto_L6115 : boolean := false;
    variable goto_L585 : boolean := false;
    variable goto_L586 : boolean := false;
    variable goto_L11 : boolean := false;
    variable goto_L13 : boolean := false;
    variable goto_L6233 : boolean := false;
    variable goto_L6266 : boolean := false;
    variable goto_L6245 : boolean := false;
    variable goto_L563 : boolean := false;
    variable goto_L0 : boolean := false;
    variable goto_L6288 : boolean := false;
    variable r6279 : std_logic_vector(0 to 513) := (others => '0');
    variable r6274 : std_logic_vector(0 to 257) := (others => '0');
    variable r6272 : std_logic_vector(0 to 1) := (others => '0');
    variable r6270 : std_logic_vector(0 to 255) := (others => '0');
    variable r6263 : std_logic_vector(0 to 513) := (others => '0');
    variable r6259 : std_logic_vector(0 to 255) := (others => '0');
    variable r6258 : std_logic_vector(0 to 257) := (others => '0');
    variable r6256 : std_logic_vector(0 to 1) := (others => '0');
    variable r6250 : std_logic_vector(0 to 5) := (others => '0');
    variable r6248 : std_logic_vector(0 to 5) := (others => '0');
    variable r6244 : std_logic_vector(0 to 255) := (others => '0');
    variable b6242 : boolean := false;
    variable b6240 : boolean := false;
    variable r6238 : std_logic_vector(0 to 511) := (others => '0');
    variable b6236 : boolean := false;
    variable r6219 : std_logic_vector(0 to 31) := (others => '0');
    variable r6215 : std_logic_vector(0 to 31) := (others => '0');
    variable r6211 : std_logic_vector(0 to 31) := (others => '0');
    variable r6207 : std_logic_vector(0 to 31) := (others => '0');
    variable r6203 : std_logic_vector(0 to 31) := (others => '0');
    variable r6199 : std_logic_vector(0 to 31) := (others => '0');
    variable r6195 : std_logic_vector(0 to 31) := (others => '0');
    variable r6191 : std_logic_vector(0 to 31) := (others => '0');
    variable r6187 : std_logic_vector(0 to 255) := (others => '0');
    variable b6184 : boolean := false;
    variable b6182 : boolean := false;
    variable b6180 : boolean := false;
    variable b6178 : boolean := false;
    variable b6176 : boolean := false;
    variable b6174 : boolean := false;
    variable b6172 : boolean := false;
    variable b6170 : boolean := false;
    variable r6168 : std_logic_vector(0 to 31) := (others => '0');
    variable r6166 : std_logic_vector(0 to 31) := (others => '0');
    variable r6164 : std_logic_vector(0 to 31) := (others => '0');
    variable r6162 : std_logic_vector(0 to 31) := (others => '0');
    variable r6160 : std_logic_vector(0 to 31) := (others => '0');
    variable r6158 : std_logic_vector(0 to 31) := (others => '0');
    variable r6156 : std_logic_vector(0 to 31) := (others => '0');
    variable r6154 : std_logic_vector(0 to 31) := (others => '0');
    variable r6150 : std_logic_vector(0 to 255) := (others => '0');
    variable b6148 : boolean := false;
    variable b6146 : boolean := false;
    variable b6144 : boolean := false;
    variable b6142 : boolean := false;
    variable b6140 : boolean := false;
    variable b6138 : boolean := false;
    variable b6136 : boolean := false;
    variable b6134 : boolean := false;
    variable r6132 : std_logic_vector(0 to 31) := (others => '0');
    variable r6130 : std_logic_vector(0 to 31) := (others => '0');
    variable r6128 : std_logic_vector(0 to 31) := (others => '0');
    variable r6126 : std_logic_vector(0 to 31) := (others => '0');
    variable r6124 : std_logic_vector(0 to 31) := (others => '0');
    variable r6122 : std_logic_vector(0 to 31) := (others => '0');
    variable r6120 : std_logic_vector(0 to 31) := (others => '0');
    variable r6118 : std_logic_vector(0 to 31) := (others => '0');
    variable r6114 : std_logic_vector(0 to 255) := (others => '0');
    variable b6112 : boolean := false;
    variable r6109 : std_logic_vector(0 to 513) := (others => '0');
    variable r6105 : std_logic_vector(0 to 255) := (others => '0');
    variable r6104 : std_logic_vector(0 to 257) := (others => '0');
    variable r6102 : std_logic_vector(0 to 1) := (others => '0');
    variable r6098 : std_logic_vector(0 to 5) := (others => '0');
    variable r6094 : std_logic_vector(0 to 255) := (others => '0');
    variable r6090 : std_logic_vector(0 to 31) := (others => '0');
    variable r1672 : std_logic_vector(0 to 5) := (others => '0');
    variable r1174 : std_logic_vector(0 to 255) := (others => '0');
    variable r1173 : std_logic_vector(0 to 31) := (others => '0');
    variable r1172 : std_logic_vector(0 to 31) := (others => '0');
    variable r1169 : std_logic_vector(0 to 255) := (others => '0');
    variable r1163 : std_logic_vector(0 to 511) := (others => '0');
    variable r660 : std_logic_vector(0 to 511) := (others => '0');
    variable b657 : boolean := false;
    variable b655 : boolean := false;
    variable b653 : boolean := false;
    variable b651 : boolean := false;
    variable b649 : boolean := false;
    variable b647 : boolean := false;
    variable b645 : boolean := false;
    variable b643 : boolean := false;
    variable b641 : boolean := false;
    variable b639 : boolean := false;
    variable b637 : boolean := false;
    variable b635 : boolean := false;
    variable b633 : boolean := false;
    variable b631 : boolean := false;
    variable b629 : boolean := false;
    variable b627 : boolean := false;
    variable r625 : std_logic_vector(0 to 31) := (others => '0');
    variable r623 : std_logic_vector(0 to 31) := (others => '0');
    variable r621 : std_logic_vector(0 to 31) := (others => '0');
    variable r619 : std_logic_vector(0 to 31) := (others => '0');
    variable r617 : std_logic_vector(0 to 31) := (others => '0');
    variable r615 : std_logic_vector(0 to 31) := (others => '0');
    variable r613 : std_logic_vector(0 to 31) := (others => '0');
    variable r611 : std_logic_vector(0 to 31) := (others => '0');
    variable r609 : std_logic_vector(0 to 31) := (others => '0');
    variable r607 : std_logic_vector(0 to 31) := (others => '0');
    variable r605 : std_logic_vector(0 to 31) := (others => '0');
    variable r603 : std_logic_vector(0 to 31) := (others => '0');
    variable r601 : std_logic_vector(0 to 31) := (others => '0');
    variable r599 : std_logic_vector(0 to 31) := (others => '0');
    variable r597 : std_logic_vector(0 to 31) := (others => '0');
    variable r595 : std_logic_vector(0 to 31) := (others => '0');
    variable r593 : std_logic_vector(0 to 31) := (others => '0');
    variable r590 : std_logic_vector(0 to 511) := (others => '0');
    variable r588 : std_logic_vector(0 to 5) := (others => '0');
    variable r584 : std_logic_vector(0 to 513) := (others => '0');
    variable r580 : std_logic_vector(0 to 255) := (others => '0');
    variable r579 : std_logic_vector(0 to 257) := (others => '0');
    variable r577 : std_logic_vector(0 to 1) := (others => '0');
    variable r571 : std_logic_vector(0 to 255) := (others => '0');
    variable r567 : std_logic_vector(0 to 5) := (others => '0');
    variable r565 : std_logic_vector(0 to 5) := (others => '0');
    variable r562 : std_logic_vector(0 to 255) := (others => '0');
    variable b22 : boolean := false;
    variable b20 : boolean := false;
    variable r18 : std_logic_vector(0 to 511) := (others => '0');
    variable b16 : boolean := false;
    variable r12 : std_logic_vector(0 to 513) := (others => '0');
    variable r10 : std_logic_vector(0 to 513) := (others => '0');
    variable r6 : std_logic_vector(0 to 255) := (others => '0');
    variable r5 : std_logic_vector(0 to 257) := (others => '0');
    variable r3 : std_logic_vector(0 to 1) := (others => '0');
    variable statevar0 : std_logic_vector(0 to 255) := (others => '0');
    variable statevar1 : std_logic_vector(0 to 511) := (others => '0');
    variable statevar2 : std_logic_vector(0 to 255) := (others => '0');
    variable statevar3 : std_logic_vector(0 to 5) := (others => '0');
    variable output_tmp : std_logic_vector(0 to 257);
  begin
    -- Read reg temps.
    control := control_flop;
    input_tmp := input_flop;
    goto_L6287 := goto_L6287_flop;
    goto_L6280 := goto_L6280_flop;
    goto_L6264 := goto_L6264_flop;
    goto_L6110 := goto_L6110_flop;
    goto_L6230 := goto_L6230_flop;
    goto_L6115 := goto_L6115_flop;
    goto_L585 := goto_L585_flop;
    goto_L586 := goto_L586_flop;
    goto_L11 := goto_L11_flop;
    goto_L13 := goto_L13_flop;
    goto_L6233 := goto_L6233_flop;
    goto_L6266 := goto_L6266_flop;
    goto_L6245 := goto_L6245_flop;
    goto_L563 := goto_L563_flop;
    goto_L0 := goto_L0_flop;
    goto_L6288 := goto_L6288_flop;
    r6279 := r6279_flop;
    r6274 := r6274_flop;
    r6272 := r6272_flop;
    r6270 := r6270_flop;
    r6263 := r6263_flop;
    r6259 := r6259_flop;
    r6258 := r6258_flop;
    r6256 := r6256_flop;
    r6250 := r6250_flop;
    r6248 := r6248_flop;
    r6244 := r6244_flop;
    b6242 := b6242_flop;
    b6240 := b6240_flop;
    r6238 := r6238_flop;
    b6236 := b6236_flop;
    r6219 := r6219_flop;
    r6215 := r6215_flop;
    r6211 := r6211_flop;
    r6207 := r6207_flop;
    r6203 := r6203_flop;
    r6199 := r6199_flop;
    r6195 := r6195_flop;
    r6191 := r6191_flop;
    r6187 := r6187_flop;
    b6184 := b6184_flop;
    b6182 := b6182_flop;
    b6180 := b6180_flop;
    b6178 := b6178_flop;
    b6176 := b6176_flop;
    b6174 := b6174_flop;
    b6172 := b6172_flop;
    b6170 := b6170_flop;
    r6168 := r6168_flop;
    r6166 := r6166_flop;
    r6164 := r6164_flop;
    r6162 := r6162_flop;
    r6160 := r6160_flop;
    r6158 := r6158_flop;
    r6156 := r6156_flop;
    r6154 := r6154_flop;
    r6150 := r6150_flop;
    b6148 := b6148_flop;
    b6146 := b6146_flop;
    b6144 := b6144_flop;
    b6142 := b6142_flop;
    b6140 := b6140_flop;
    b6138 := b6138_flop;
    b6136 := b6136_flop;
    b6134 := b6134_flop;
    r6132 := r6132_flop;
    r6130 := r6130_flop;
    r6128 := r6128_flop;
    r6126 := r6126_flop;
    r6124 := r6124_flop;
    r6122 := r6122_flop;
    r6120 := r6120_flop;
    r6118 := r6118_flop;
    r6114 := r6114_flop;
    b6112 := b6112_flop;
    r6109 := r6109_flop;
    r6105 := r6105_flop;
    r6104 := r6104_flop;
    r6102 := r6102_flop;
    r6098 := r6098_flop;
    r6094 := r6094_flop;
    r6090 := r6090_flop;
    r1672 := r1672_flop;
    r1174 := r1174_flop;
    r1173 := r1173_flop;
    r1172 := r1172_flop;
    r1169 := r1169_flop;
    r1163 := r1163_flop;
    r660 := r660_flop;
    b657 := b657_flop;
    b655 := b655_flop;
    b653 := b653_flop;
    b651 := b651_flop;
    b649 := b649_flop;
    b647 := b647_flop;
    b645 := b645_flop;
    b643 := b643_flop;
    b641 := b641_flop;
    b639 := b639_flop;
    b637 := b637_flop;
    b635 := b635_flop;
    b633 := b633_flop;
    b631 := b631_flop;
    b629 := b629_flop;
    b627 := b627_flop;
    r625 := r625_flop;
    r623 := r623_flop;
    r621 := r621_flop;
    r619 := r619_flop;
    r617 := r617_flop;
    r615 := r615_flop;
    r613 := r613_flop;
    r611 := r611_flop;
    r609 := r609_flop;
    r607 := r607_flop;
    r605 := r605_flop;
    r603 := r603_flop;
    r601 := r601_flop;
    r599 := r599_flop;
    r597 := r597_flop;
    r595 := r595_flop;
    r593 := r593_flop;
    r590 := r590_flop;
    r588 := r588_flop;
    r584 := r584_flop;
    r580 := r580_flop;
    r579 := r579_flop;
    r577 := r577_flop;
    r571 := r571_flop;
    r567 := r567_flop;
    r565 := r565_flop;
    r562 := r562_flop;
    b22 := b22_flop;
    b20 := b20_flop;
    r18 := r18_flop;
    b16 := b16_flop;
    r12 := r12_flop;
    r10 := r10_flop;
    r6 := r6_flop;
    r5 := r5_flop;
    r3 := r3_flop;
    statevar0 := statevar0_flop;
    statevar1 := statevar1_flop;
    statevar2 := statevar2_flop;
    statevar3 := statevar3_flop;
    output_tmp := (others => '0');
    -- Loop body.
    goto_L6287 := false;
    goto_L6280 := false;
    goto_L6264 := false;
    goto_L6110 := false;
    goto_L6230 := false;
    goto_L6115 := false;
    goto_L585 := false;
    goto_L586 := false;
    goto_L11 := false;
    goto_L13 := false;
    goto_L6233 := false;
    goto_L6266 := false;
    goto_L6245 := false;
    goto_L563 := false;
    goto_L0 := false;
    goto_L6288 := false;
    null; -- label L6287
    -- ENTER
    goto_L0 := (control = STATE0);
    if (NOT goto_L0) then
      goto_L11 := (control = STATE11);
      if (NOT goto_L11) then
        goto_L585 := (control = STATE585);
        if (NOT goto_L585) then
          goto_L6110 := (control = STATE6110);
          if (NOT goto_L6110) then
            goto_L6264 := (control = STATE6264);
            if (NOT goto_L6264) then
              goto_L6280 := (control = STATE6280);
              null; -- label L6280
              r6279 := input_tmp;
              -- got i@1V4 in r6279
              r12 := r6279;
              goto_L13 := true;
            end if;
            goto_L13 := goto_L13;
            if (NOT goto_L13) then
              null; -- label L6264
              r6263 := input_tmp;
              goto_L586 := true;
            end if;
            goto_L586 := goto_L586;
          end if;
          goto_L586 := goto_L586;
          if (NOT goto_L586) then
            goto_L13 := goto_L13;
            if (NOT goto_L13) then
              null; -- label L6110
              r6109 := input_tmp;
              -- got ctr@1VS in r588
              b6112 := ("111111" = r588(0 to 5));
              goto_L6115 := b6112;
              if (NOT goto_L6115) then
                goto_L6230 := (NOT b6112);
                null; -- label L6230
                -- alt exit (no match)
                goto_L586 := true;
              end if;
              goto_L586 := goto_L586;
              if (NOT goto_L586) then
                null; -- label L6115
                r6114 := statevar2;
                -- got $19@1VU in r6114
                -- final pat
                r6118 := r6114(0 to 31);
                r6120 := r6114(32 to 63);
                r6122 := r6114(64 to 95);
                r6124 := r6114(96 to 127);
                r6126 := r6114(128 to 159);
                r6128 := r6114(160 to 191);
                r6130 := r6114(192 to 223);
                r6132 := r6114(224 to 255);
                b6134 := true;
                b6136 := true;
                b6138 := true;
                b6140 := true;
                b6142 := true;
                b6144 := true;
                b6146 := true;
                b6148 := true;
                r6150 := statevar0;
                -- got $18@207 in r6150
                -- final pat
                r6154 := r6150(0 to 31);
                r6156 := r6150(32 to 63);
                r6158 := r6150(64 to 95);
                r6160 := r6150(96 to 127);
                r6162 := r6150(128 to 159);
                r6164 := r6150(160 to 191);
                r6166 := r6150(192 to 223);
                r6168 := r6150(224 to 255);
                b6170 := true;
                b6172 := true;
                b6174 := true;
                b6176 := true;
                b6178 := true;
                b6180 := true;
                b6182 := true;
                b6184 := true;
                null;
                null;
                -- got a@208 in r6154
                -- got h1@1VV in r6118
                r6191 := w32Plus(r6154,r6118);
                -- got b@209 in r6156
                -- got h2@200 in r6120
                r6195 := w32Plus(r6156,r6120);
                -- got c@20A in r6158
                -- got h3@201 in r6122
                r6199 := w32Plus(r6158,r6122);
                -- got d@20B in r6160
                -- got h4@202 in r6124
                r6203 := w32Plus(r6160,r6124);
                -- got e@20C in r6162
                -- got h5@203 in r6126
                r6207 := w32Plus(r6162,r6126);
                -- got f@20D in r6164
                -- got h6@204 in r6128
                r6211 := w32Plus(r6164,r6128);
                -- got g@20E in r6166
                -- got h7@205 in r6130
                r6215 := w32Plus(r6166,r6130);
                -- got h@20F in r6168
                -- got h8@206 in r6132
                r6219 := w32Plus(r6168,r6132);
                r6187 := (r6191 & r6195 & r6199 & r6203 & r6207 & r6211 & r6215 & r6219);
                statevar2 := r6187;
                null;
                -- end case
                null;
                -- end case
                -- got i@1VT in r6109
                r12 := r6109;
                goto_L13 := true;
              end if;
              goto_L13 := goto_L13;
            end if;
            goto_L13 := goto_L13;
            if (NOT goto_L13) then
              goto_L586 := goto_L586;
            end if;
            goto_L586 := goto_L586;
          end if;
          goto_L586 := goto_L586;
          if (NOT goto_L586) then
            goto_L13 := goto_L13;
          end if;
          goto_L13 := goto_L13;
        end if;
        goto_L13 := goto_L13;
        if (NOT goto_L13) then
          goto_L586 := goto_L586;
          if (NOT goto_L586) then
            null; -- label L585
            r584 := input_tmp;
            goto_L586 := true;
          end if;
          goto_L586 := goto_L586;
          null; -- label L586
          -- Main.loop in
          r588 := statevar3;
          r590 := statevar1;
          -- got s@1V6 in r590
          -- final pat
          r595 := r590(0 to 31);
          r597 := r590(32 to 63);
          r599 := r590(64 to 95);
          r601 := r590(96 to 127);
          r603 := r590(128 to 159);
          r605 := r590(160 to 191);
          r607 := r590(192 to 223);
          r609 := r590(224 to 255);
          r611 := r590(256 to 287);
          r613 := r590(288 to 319);
          r615 := r590(320 to 351);
          r617 := r590(352 to 383);
          r619 := r590(384 to 415);
          r621 := r590(416 to 447);
          r623 := r590(448 to 479);
          r625 := r590(480 to 511);
          b627 := true;
          b629 := true;
          b631 := true;
          b633 := true;
          b635 := true;
          b637 := true;
          b639 := true;
          b641 := true;
          b643 := true;
          b645 := true;
          b647 := true;
          b649 := true;
          b651 := true;
          b653 := true;
          b655 := true;
          b657 := true;
          -- got s@1V6 in r590
          r1163 := rewire_Main.updateSched_659(r590);
          statevar1 := r1163;
          -- got w00@1V7 in r595
          r593 := r595;
          -- end case
          r1169 := statevar0;
          -- got ctr@1V5 in r588
          r6090 := rewire_Main.seed_1671(r588);
          -- got $12@1VO in r593
          -- got s@1VP in r1169
          r6094 := rewire_Main.step256_1171(r6090,r593,r1169);
          statevar0 := r6094;
          -- got ctr@1V5 in r588
          r6098 := incCtr(r588);
          statevar3 := r6098;
          -- got ctr@1V5 in r588
          r6102 := "10";
          r6105 := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
          r6104 := (r6102 & r6105);
          output_tmp := r6104;
          control := STATE6110;
          goto_L6288 := true;
        end if;
        goto_L6288 := goto_L6288;
      end if;
      goto_L6288 := goto_L6288;
      if (NOT goto_L6288) then
        goto_L13 := goto_L13;
        if (NOT goto_L13) then
          null; -- label L11
          r10 := input_tmp;
          -- got i@1UK in r10
          r12 := r10;
          goto_L13 := true;
        end if;
        goto_L13 := goto_L13;
        null; -- label L13
        -- Main.dev in
        -- got $16@1UL in r12
        b16 := ("00" = r12(0 to 1));
        r18 := r12(2 to 513);
        b20 := true;
        b22 := (b16 AND b20);
        goto_L563 := b22;
        if (NOT goto_L563) then
          goto_L6233 := (NOT b22);
          null; -- label L6233
          -- alt exit (no match)
          -- got $16@1UL in r12
          b6236 := ("01" = r12(0 to 1));
          r6238 := r12(2 to 513);
          b6240 := true;
          b6242 := (b6236 AND b6240);
          goto_L6245 := b6242;
          if (NOT goto_L6245) then
            goto_L6266 := (NOT b6242);
            null; -- label L6266
            -- alt exit (no match)
            -- got $16@1UL in r12
            -- final pat
            r6270 := statevar2;
            r6272 := "00";
            null;
            -- got h_n@1V3 in r6270
            r6274 := (r6272 & r6270);
            output_tmp := r6274;
            control := STATE6280;
            goto_L6288 := true;
          end if;
          goto_L6288 := goto_L6288;
          if (NOT goto_L6288) then
            null; -- label L6245
            r6244 := statevar2;
            -- got hi_1@1UU in r6244
            statevar0 := r6244;
            r6248 := "000000";
            null;
            r6250 := (r6248);
            statevar3 := r6250;
            -- got hw32@1UT in r6238
            statevar1 := r6238;
            r6256 := "01";
            r6259 := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
            r6258 := (r6256 & r6259);
            output_tmp := r6258;
            control := STATE6264;
            goto_L6288 := true;
          end if;
          goto_L6288 := goto_L6288;
        end if;
        goto_L6288 := goto_L6288;
        if (NOT goto_L6288) then
          null; -- label L563
          r562 := rewire_Main.initialSHA256State_24;
          statevar2 := r562;
          r565 := "000000";
          null;
          r567 := (r565);
          statevar3 := r567;
          r571 := statevar2;
          -- got hi_1@1UP in r571
          statevar0 := r571;
          -- got hw32@1UM in r18
          statevar1 := r18;
          r577 := "01";
          r580 := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
          r579 := (r577 & r580);
          output_tmp := r579;
          control := STATE585;
          goto_L6288 := true;
        end if;
        goto_L6288 := goto_L6288;
      end if;
      goto_L6288 := goto_L6288;
    end if;
    goto_L6288 := goto_L6288;
    if (NOT goto_L6288) then
      null; -- label L0
      -- START
      -- Main.devsha256' in
      r3 := "01";
      r6 := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      r5 := (r3 & r6);
      output_tmp := r5;
      control := STATE11;
      goto_L6288 := true;
    end if;
    goto_L6288 := goto_L6288;
    null; -- label L6288
    -- EXIT
    -- Write back reg temps.
    control_flop_next <= control;
    goto_L6287_flop_next <= goto_L6287;
    goto_L6280_flop_next <= goto_L6280;
    goto_L6264_flop_next <= goto_L6264;
    goto_L6110_flop_next <= goto_L6110;
    goto_L6230_flop_next <= goto_L6230;
    goto_L6115_flop_next <= goto_L6115;
    goto_L585_flop_next <= goto_L585;
    goto_L586_flop_next <= goto_L586;
    goto_L11_flop_next <= goto_L11;
    goto_L13_flop_next <= goto_L13;
    goto_L6233_flop_next <= goto_L6233;
    goto_L6266_flop_next <= goto_L6266;
    goto_L6245_flop_next <= goto_L6245;
    goto_L563_flop_next <= goto_L563;
    goto_L0_flop_next <= goto_L0;
    goto_L6288_flop_next <= goto_L6288;
    r6279_flop_next <= r6279;
    r6274_flop_next <= r6274;
    r6272_flop_next <= r6272;
    r6270_flop_next <= r6270;
    r6263_flop_next <= r6263;
    r6259_flop_next <= r6259;
    r6258_flop_next <= r6258;
    r6256_flop_next <= r6256;
    r6250_flop_next <= r6250;
    r6248_flop_next <= r6248;
    r6244_flop_next <= r6244;
    b6242_flop_next <= b6242;
    b6240_flop_next <= b6240;
    r6238_flop_next <= r6238;
    b6236_flop_next <= b6236;
    r6219_flop_next <= r6219;
    r6215_flop_next <= r6215;
    r6211_flop_next <= r6211;
    r6207_flop_next <= r6207;
    r6203_flop_next <= r6203;
    r6199_flop_next <= r6199;
    r6195_flop_next <= r6195;
    r6191_flop_next <= r6191;
    r6187_flop_next <= r6187;
    b6184_flop_next <= b6184;
    b6182_flop_next <= b6182;
    b6180_flop_next <= b6180;
    b6178_flop_next <= b6178;
    b6176_flop_next <= b6176;
    b6174_flop_next <= b6174;
    b6172_flop_next <= b6172;
    b6170_flop_next <= b6170;
    r6168_flop_next <= r6168;
    r6166_flop_next <= r6166;
    r6164_flop_next <= r6164;
    r6162_flop_next <= r6162;
    r6160_flop_next <= r6160;
    r6158_flop_next <= r6158;
    r6156_flop_next <= r6156;
    r6154_flop_next <= r6154;
    r6150_flop_next <= r6150;
    b6148_flop_next <= b6148;
    b6146_flop_next <= b6146;
    b6144_flop_next <= b6144;
    b6142_flop_next <= b6142;
    b6140_flop_next <= b6140;
    b6138_flop_next <= b6138;
    b6136_flop_next <= b6136;
    b6134_flop_next <= b6134;
    r6132_flop_next <= r6132;
    r6130_flop_next <= r6130;
    r6128_flop_next <= r6128;
    r6126_flop_next <= r6126;
    r6124_flop_next <= r6124;
    r6122_flop_next <= r6122;
    r6120_flop_next <= r6120;
    r6118_flop_next <= r6118;
    r6114_flop_next <= r6114;
    b6112_flop_next <= b6112;
    r6109_flop_next <= r6109;
    r6105_flop_next <= r6105;
    r6104_flop_next <= r6104;
    r6102_flop_next <= r6102;
    r6098_flop_next <= r6098;
    r6094_flop_next <= r6094;
    r6090_flop_next <= r6090;
    r1672_flop_next <= r1672;
    r1174_flop_next <= r1174;
    r1173_flop_next <= r1173;
    r1172_flop_next <= r1172;
    r1169_flop_next <= r1169;
    r1163_flop_next <= r1163;
    r660_flop_next <= r660;
    b657_flop_next <= b657;
    b655_flop_next <= b655;
    b653_flop_next <= b653;
    b651_flop_next <= b651;
    b649_flop_next <= b649;
    b647_flop_next <= b647;
    b645_flop_next <= b645;
    b643_flop_next <= b643;
    b641_flop_next <= b641;
    b639_flop_next <= b639;
    b637_flop_next <= b637;
    b635_flop_next <= b635;
    b633_flop_next <= b633;
    b631_flop_next <= b631;
    b629_flop_next <= b629;
    b627_flop_next <= b627;
    r625_flop_next <= r625;
    r623_flop_next <= r623;
    r621_flop_next <= r621;
    r619_flop_next <= r619;
    r617_flop_next <= r617;
    r615_flop_next <= r615;
    r613_flop_next <= r613;
    r611_flop_next <= r611;
    r609_flop_next <= r609;
    r607_flop_next <= r607;
    r605_flop_next <= r605;
    r603_flop_next <= r603;
    r601_flop_next <= r601;
    r599_flop_next <= r599;
    r597_flop_next <= r597;
    r595_flop_next <= r595;
    r593_flop_next <= r593;
    r590_flop_next <= r590;
    r588_flop_next <= r588;
    r584_flop_next <= r584;
    r580_flop_next <= r580;
    r579_flop_next <= r579;
    r577_flop_next <= r577;
    r571_flop_next <= r571;
    r567_flop_next <= r567;
    r565_flop_next <= r565;
    r562_flop_next <= r562;
    b22_flop_next <= b22;
    b20_flop_next <= b20;
    r18_flop_next <= r18;
    b16_flop_next <= b16;
    r12_flop_next <= r12;
    r10_flop_next <= r10;
    r6_flop_next <= r6;
    r5_flop_next <= r5;
    r3_flop_next <= r3;
    statevar0_flop_next <= statevar0;
    statevar1_flop_next <= statevar1;
    statevar2_flop_next <= statevar2;
    statevar3_flop_next <= statevar3;
    -- Update output line.
    output <= output_tmp;
  end process;

  -- Flip flop update process.
  process (clk,input,goto_L6287_flop_next,goto_L6280_flop_next,goto_L6264_flop_next,goto_L6110_flop_next,goto_L6230_flop_next,goto_L6115_flop_next,goto_L585_flop_next,goto_L586_flop_next,goto_L11_flop_next,goto_L13_flop_next,goto_L6233_flop_next,goto_L6266_flop_next,goto_L6245_flop_next,goto_L563_flop_next,goto_L0_flop_next,goto_L6288_flop_next,r6279_flop_next,r6274_flop_next,r6272_flop_next,r6270_flop_next,r6263_flop_next,r6259_flop_next,r6258_flop_next,r6256_flop_next,r6250_flop_next,r6248_flop_next,r6244_flop_next,b6242_flop_next,b6240_flop_next,r6238_flop_next,b6236_flop_next,r6219_flop_next,r6215_flop_next,r6211_flop_next,r6207_flop_next,r6203_flop_next,r6199_flop_next,r6195_flop_next,r6191_flop_next,r6187_flop_next,b6184_flop_next,b6182_flop_next,b6180_flop_next,b6178_flop_next,b6176_flop_next,b6174_flop_next,b6172_flop_next,b6170_flop_next,r6168_flop_next,r6166_flop_next,r6164_flop_next,r6162_flop_next,r6160_flop_next,r6158_flop_next,r6156_flop_next,r6154_flop_next,r6150_flop_next,b6148_flop_next,b6146_flop_next,b6144_flop_next,b6142_flop_next,b6140_flop_next,b6138_flop_next,b6136_flop_next,b6134_flop_next,r6132_flop_next,r6130_flop_next,r6128_flop_next,r6126_flop_next,r6124_flop_next,r6122_flop_next,r6120_flop_next,r6118_flop_next,r6114_flop_next,b6112_flop_next,r6109_flop_next,r6105_flop_next,r6104_flop_next,r6102_flop_next,r6098_flop_next,r6094_flop_next,r6090_flop_next,r1672_flop_next,r1174_flop_next,r1173_flop_next,r1172_flop_next,r1169_flop_next,r1163_flop_next,r660_flop_next,b657_flop_next,b655_flop_next,b653_flop_next,b651_flop_next,b649_flop_next,b647_flop_next,b645_flop_next,b643_flop_next,b641_flop_next,b639_flop_next,b637_flop_next,b635_flop_next,b633_flop_next,b631_flop_next,b629_flop_next,b627_flop_next,r625_flop_next,r623_flop_next,r621_flop_next,r619_flop_next,r617_flop_next,r615_flop_next,r613_flop_next,r611_flop_next,r609_flop_next,r607_flop_next,r605_flop_next,r603_flop_next,r601_flop_next,r599_flop_next,r597_flop_next,r595_flop_next,r593_flop_next,r590_flop_next,r588_flop_next,r584_flop_next,r580_flop_next,r579_flop_next,r577_flop_next,r571_flop_next,r567_flop_next,r565_flop_next,r562_flop_next,b22_flop_next,b20_flop_next,r18_flop_next,b16_flop_next,r12_flop_next,r10_flop_next,r6_flop_next,r5_flop_next,r3_flop_next,statevar0_flop_next,statevar1_flop_next,statevar2_flop_next,statevar3_flop_next)
  begin
    if clk'event and clk='1' then
      input_flop <= input;
      control_flop <= control_flop_next;
      goto_L6287_flop <= goto_L6287_flop_next;
      goto_L6280_flop <= goto_L6280_flop_next;
      goto_L6264_flop <= goto_L6264_flop_next;
      goto_L6110_flop <= goto_L6110_flop_next;
      goto_L6230_flop <= goto_L6230_flop_next;
      goto_L6115_flop <= goto_L6115_flop_next;
      goto_L585_flop <= goto_L585_flop_next;
      goto_L586_flop <= goto_L586_flop_next;
      goto_L11_flop <= goto_L11_flop_next;
      goto_L13_flop <= goto_L13_flop_next;
      goto_L6233_flop <= goto_L6233_flop_next;
      goto_L6266_flop <= goto_L6266_flop_next;
      goto_L6245_flop <= goto_L6245_flop_next;
      goto_L563_flop <= goto_L563_flop_next;
      goto_L0_flop <= goto_L0_flop_next;
      goto_L6288_flop <= goto_L6288_flop_next;
      r6279_flop <= r6279_flop_next;
      r6274_flop <= r6274_flop_next;
      r6272_flop <= r6272_flop_next;
      r6270_flop <= r6270_flop_next;
      r6263_flop <= r6263_flop_next;
      r6259_flop <= r6259_flop_next;
      r6258_flop <= r6258_flop_next;
      r6256_flop <= r6256_flop_next;
      r6250_flop <= r6250_flop_next;
      r6248_flop <= r6248_flop_next;
      r6244_flop <= r6244_flop_next;
      b6242_flop <= b6242_flop_next;
      b6240_flop <= b6240_flop_next;
      r6238_flop <= r6238_flop_next;
      b6236_flop <= b6236_flop_next;
      r6219_flop <= r6219_flop_next;
      r6215_flop <= r6215_flop_next;
      r6211_flop <= r6211_flop_next;
      r6207_flop <= r6207_flop_next;
      r6203_flop <= r6203_flop_next;
      r6199_flop <= r6199_flop_next;
      r6195_flop <= r6195_flop_next;
      r6191_flop <= r6191_flop_next;
      r6187_flop <= r6187_flop_next;
      b6184_flop <= b6184_flop_next;
      b6182_flop <= b6182_flop_next;
      b6180_flop <= b6180_flop_next;
      b6178_flop <= b6178_flop_next;
      b6176_flop <= b6176_flop_next;
      b6174_flop <= b6174_flop_next;
      b6172_flop <= b6172_flop_next;
      b6170_flop <= b6170_flop_next;
      r6168_flop <= r6168_flop_next;
      r6166_flop <= r6166_flop_next;
      r6164_flop <= r6164_flop_next;
      r6162_flop <= r6162_flop_next;
      r6160_flop <= r6160_flop_next;
      r6158_flop <= r6158_flop_next;
      r6156_flop <= r6156_flop_next;
      r6154_flop <= r6154_flop_next;
      r6150_flop <= r6150_flop_next;
      b6148_flop <= b6148_flop_next;
      b6146_flop <= b6146_flop_next;
      b6144_flop <= b6144_flop_next;
      b6142_flop <= b6142_flop_next;
      b6140_flop <= b6140_flop_next;
      b6138_flop <= b6138_flop_next;
      b6136_flop <= b6136_flop_next;
      b6134_flop <= b6134_flop_next;
      r6132_flop <= r6132_flop_next;
      r6130_flop <= r6130_flop_next;
      r6128_flop <= r6128_flop_next;
      r6126_flop <= r6126_flop_next;
      r6124_flop <= r6124_flop_next;
      r6122_flop <= r6122_flop_next;
      r6120_flop <= r6120_flop_next;
      r6118_flop <= r6118_flop_next;
      r6114_flop <= r6114_flop_next;
      b6112_flop <= b6112_flop_next;
      r6109_flop <= r6109_flop_next;
      r6105_flop <= r6105_flop_next;
      r6104_flop <= r6104_flop_next;
      r6102_flop <= r6102_flop_next;
      r6098_flop <= r6098_flop_next;
      r6094_flop <= r6094_flop_next;
      r6090_flop <= r6090_flop_next;
      r1672_flop <= r1672_flop_next;
      r1174_flop <= r1174_flop_next;
      r1173_flop <= r1173_flop_next;
      r1172_flop <= r1172_flop_next;
      r1169_flop <= r1169_flop_next;
      r1163_flop <= r1163_flop_next;
      r660_flop <= r660_flop_next;
      b657_flop <= b657_flop_next;
      b655_flop <= b655_flop_next;
      b653_flop <= b653_flop_next;
      b651_flop <= b651_flop_next;
      b649_flop <= b649_flop_next;
      b647_flop <= b647_flop_next;
      b645_flop <= b645_flop_next;
      b643_flop <= b643_flop_next;
      b641_flop <= b641_flop_next;
      b639_flop <= b639_flop_next;
      b637_flop <= b637_flop_next;
      b635_flop <= b635_flop_next;
      b633_flop <= b633_flop_next;
      b631_flop <= b631_flop_next;
      b629_flop <= b629_flop_next;
      b627_flop <= b627_flop_next;
      r625_flop <= r625_flop_next;
      r623_flop <= r623_flop_next;
      r621_flop <= r621_flop_next;
      r619_flop <= r619_flop_next;
      r617_flop <= r617_flop_next;
      r615_flop <= r615_flop_next;
      r613_flop <= r613_flop_next;
      r611_flop <= r611_flop_next;
      r609_flop <= r609_flop_next;
      r607_flop <= r607_flop_next;
      r605_flop <= r605_flop_next;
      r603_flop <= r603_flop_next;
      r601_flop <= r601_flop_next;
      r599_flop <= r599_flop_next;
      r597_flop <= r597_flop_next;
      r595_flop <= r595_flop_next;
      r593_flop <= r593_flop_next;
      r590_flop <= r590_flop_next;
      r588_flop <= r588_flop_next;
      r584_flop <= r584_flop_next;
      r580_flop <= r580_flop_next;
      r579_flop <= r579_flop_next;
      r577_flop <= r577_flop_next;
      r571_flop <= r571_flop_next;
      r567_flop <= r567_flop_next;
      r565_flop <= r565_flop_next;
      r562_flop <= r562_flop_next;
      b22_flop <= b22_flop_next;
      b20_flop <= b20_flop_next;
      r18_flop <= r18_flop_next;
      b16_flop <= b16_flop_next;
      r12_flop <= r12_flop_next;
      r10_flop <= r10_flop_next;
      r6_flop <= r6_flop_next;
      r5_flop <= r5_flop_next;
      r3_flop <= r3_flop_next;
      statevar0_flop <= statevar0_flop_next;
      statevar1_flop <= statevar1_flop_next;
      statevar2_flop <= statevar2_flop_next;
      statevar3_flop <= statevar3_flop_next;
    end if;
  end process;

end behavioral;
