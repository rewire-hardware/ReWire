library ieee;
use ieee.std_logic_1164.all;
-- Comment out the following line if VHDL primitives are not in use.
use work.prims.all;
entity rewire is
  Port ( clk : in std_logic ;
         input : in std_logic_vector (0 to 52);
         output : out std_logic_vector (0 to 36));
end rewire;

architecture behavioral of rewire is
  type control_state is (STATE0,STATE11,STATE581,STATE597);
  function rewire_Maincrossbar_32(r33 : std_logic_vector ; r34 : std_logic_vector) return std_logic_vector;
  function rewire_Maincrossbar_32(r33 : std_logic_vector ; r34 : std_logic_vector) return std_logic_vector
  is
    variable r573 : std_logic_vector(0 to 35) := (others => '0');
    variable b572 : boolean := false;
    variable b571 : boolean := false;
    variable b570 : boolean := false;
    variable r569 : std_logic_vector(0 to 8) := (others => '0');
    variable r568 : std_logic_vector(0 to 8) := (others => '0');
    variable b567 : boolean := false;
    variable r566 : std_logic_vector(0 to 35) := (others => '0');
    variable r565 : std_logic_vector(0 to 17) := (others => '0');
    variable b564 : boolean := false;
    variable b563 : boolean := false;
    variable b562 : boolean := false;
    variable b561 : boolean := false;
    variable r560 : std_logic_vector(0 to 0) := (others => '0');
    variable r559 : std_logic_vector(0 to 8) := (others => '0');
    variable r558 : std_logic_vector(0 to 8) := (others => '0');
    variable b557 : boolean := false;
    variable r556 : std_logic_vector(0 to 17) := (others => '0');
    variable r555 : std_logic_vector(0 to 18) := (others => '0');
    variable r554 : std_logic_vector(0 to 17) := (others => '0');
    variable b553 : boolean := false;
    variable b552 : boolean := false;
    variable b551 : boolean := false;
    variable b550 : boolean := false;
    variable r549 : std_logic_vector(0 to 0) := (others => '0');
    variable r548 : std_logic_vector(0 to 8) := (others => '0');
    variable r547 : std_logic_vector(0 to 8) := (others => '0');
    variable b546 : boolean := false;
    variable r545 : std_logic_vector(0 to 17) := (others => '0');
    variable r544 : std_logic_vector(0 to 18) := (others => '0');
    variable b543 : boolean := false;
    variable b542 : boolean := false;
    variable b541 : boolean := false;
    variable r540 : std_logic_vector(0 to 8) := (others => '0');
    variable r539 : std_logic_vector(0 to 8) := (others => '0');
    variable b538 : boolean := false;
    variable r537 : std_logic_vector(0 to 35) := (others => '0');
    variable r536 : std_logic_vector(0 to 17) := (others => '0');
    variable b535 : boolean := false;
    variable b534 : boolean := false;
    variable b533 : boolean := false;
    variable b532 : boolean := false;
    variable r531 : std_logic_vector(0 to 0) := (others => '0');
    variable r530 : std_logic_vector(0 to 8) := (others => '0');
    variable r529 : std_logic_vector(0 to 8) := (others => '0');
    variable b528 : boolean := false;
    variable r527 : std_logic_vector(0 to 17) := (others => '0');
    variable r526 : std_logic_vector(0 to 18) := (others => '0');
    variable r525 : std_logic_vector(0 to 17) := (others => '0');
    variable b524 : boolean := false;
    variable b523 : boolean := false;
    variable b522 : boolean := false;
    variable b521 : boolean := false;
    variable r520 : std_logic_vector(0 to 0) := (others => '0');
    variable r519 : std_logic_vector(0 to 8) := (others => '0');
    variable r518 : std_logic_vector(0 to 8) := (others => '0');
    variable b517 : boolean := false;
    variable r516 : std_logic_vector(0 to 17) := (others => '0');
    variable r515 : std_logic_vector(0 to 18) := (others => '0');
    variable b514 : boolean := false;
    variable b513 : boolean := false;
    variable b512 : boolean := false;
    variable r511 : std_logic_vector(0 to 8) := (others => '0');
    variable r510 : std_logic_vector(0 to 8) := (others => '0');
    variable b509 : boolean := false;
    variable r508 : std_logic_vector(0 to 35) := (others => '0');
    variable r507 : std_logic_vector(0 to 17) := (others => '0');
    variable b506 : boolean := false;
    variable b505 : boolean := false;
    variable b504 : boolean := false;
    variable b503 : boolean := false;
    variable r502 : std_logic_vector(0 to 0) := (others => '0');
    variable r501 : std_logic_vector(0 to 8) := (others => '0');
    variable r500 : std_logic_vector(0 to 8) := (others => '0');
    variable b499 : boolean := false;
    variable r498 : std_logic_vector(0 to 17) := (others => '0');
    variable r497 : std_logic_vector(0 to 18) := (others => '0');
    variable r496 : std_logic_vector(0 to 17) := (others => '0');
    variable b495 : boolean := false;
    variable b494 : boolean := false;
    variable b493 : boolean := false;
    variable b492 : boolean := false;
    variable r491 : std_logic_vector(0 to 0) := (others => '0');
    variable r490 : std_logic_vector(0 to 8) := (others => '0');
    variable r489 : std_logic_vector(0 to 8) := (others => '0');
    variable b488 : boolean := false;
    variable r487 : std_logic_vector(0 to 17) := (others => '0');
    variable r486 : std_logic_vector(0 to 18) := (others => '0');
    variable b485 : boolean := false;
    variable b484 : boolean := false;
    variable b483 : boolean := false;
    variable r482 : std_logic_vector(0 to 8) := (others => '0');
    variable r481 : std_logic_vector(0 to 8) := (others => '0');
    variable b480 : boolean := false;
    variable r479 : std_logic_vector(0 to 35) := (others => '0');
    variable r478 : std_logic_vector(0 to 17) := (others => '0');
    variable b477 : boolean := false;
    variable b476 : boolean := false;
    variable b475 : boolean := false;
    variable b474 : boolean := false;
    variable r473 : std_logic_vector(0 to 0) := (others => '0');
    variable r472 : std_logic_vector(0 to 8) := (others => '0');
    variable r471 : std_logic_vector(0 to 8) := (others => '0');
    variable b470 : boolean := false;
    variable r469 : std_logic_vector(0 to 17) := (others => '0');
    variable r468 : std_logic_vector(0 to 7) := (others => '0');
    variable r467 : std_logic_vector(0 to 8) := (others => '0');
    variable r466 : std_logic_vector(0 to 0) := (others => '0');
    variable r465 : std_logic_vector(0 to 18) := (others => '0');
    variable r464 : std_logic_vector(0 to 17) := (others => '0');
    variable b463 : boolean := false;
    variable b462 : boolean := false;
    variable b461 : boolean := false;
    variable b460 : boolean := false;
    variable r459 : std_logic_vector(0 to 0) := (others => '0');
    variable r458 : std_logic_vector(0 to 8) := (others => '0');
    variable r457 : std_logic_vector(0 to 8) := (others => '0');
    variable b456 : boolean := false;
    variable r455 : std_logic_vector(0 to 17) := (others => '0');
    variable r454 : std_logic_vector(0 to 7) := (others => '0');
    variable r453 : std_logic_vector(0 to 8) := (others => '0');
    variable r452 : std_logic_vector(0 to 0) := (others => '0');
    variable r451 : std_logic_vector(0 to 18) := (others => '0');
    variable b450 : boolean := false;
    variable b449 : boolean := false;
    variable b448 : boolean := false;
    variable r447 : std_logic_vector(0 to 8) := (others => '0');
    variable r446 : std_logic_vector(0 to 8) := (others => '0');
    variable b445 : boolean := false;
    variable r444 : std_logic_vector(0 to 35) := (others => '0');
    variable r443 : std_logic_vector(0 to 17) := (others => '0');
    variable b442 : boolean := false;
    variable b441 : boolean := false;
    variable b440 : boolean := false;
    variable b439 : boolean := false;
    variable r438 : std_logic_vector(0 to 0) := (others => '0');
    variable r437 : std_logic_vector(0 to 8) := (others => '0');
    variable r436 : std_logic_vector(0 to 8) := (others => '0');
    variable b435 : boolean := false;
    variable r434 : std_logic_vector(0 to 17) := (others => '0');
    variable r433 : std_logic_vector(0 to 18) := (others => '0');
    variable r432 : std_logic_vector(0 to 17) := (others => '0');
    variable b431 : boolean := false;
    variable b430 : boolean := false;
    variable b429 : boolean := false;
    variable b428 : boolean := false;
    variable r427 : std_logic_vector(0 to 0) := (others => '0');
    variable r426 : std_logic_vector(0 to 8) := (others => '0');
    variable r425 : std_logic_vector(0 to 8) := (others => '0');
    variable b424 : boolean := false;
    variable r423 : std_logic_vector(0 to 17) := (others => '0');
    variable r422 : std_logic_vector(0 to 18) := (others => '0');
    variable b421 : boolean := false;
    variable b420 : boolean := false;
    variable b419 : boolean := false;
    variable r418 : std_logic_vector(0 to 8) := (others => '0');
    variable r417 : std_logic_vector(0 to 8) := (others => '0');
    variable b416 : boolean := false;
    variable r415 : std_logic_vector(0 to 35) := (others => '0');
    variable r414 : std_logic_vector(0 to 17) := (others => '0');
    variable b413 : boolean := false;
    variable b412 : boolean := false;
    variable b411 : boolean := false;
    variable b410 : boolean := false;
    variable r409 : std_logic_vector(0 to 0) := (others => '0');
    variable r408 : std_logic_vector(0 to 8) := (others => '0');
    variable r407 : std_logic_vector(0 to 8) := (others => '0');
    variable b406 : boolean := false;
    variable r405 : std_logic_vector(0 to 17) := (others => '0');
    variable r404 : std_logic_vector(0 to 18) := (others => '0');
    variable r403 : std_logic_vector(0 to 17) := (others => '0');
    variable b402 : boolean := false;
    variable b401 : boolean := false;
    variable b400 : boolean := false;
    variable b399 : boolean := false;
    variable r398 : std_logic_vector(0 to 0) := (others => '0');
    variable r397 : std_logic_vector(0 to 8) := (others => '0');
    variable r396 : std_logic_vector(0 to 8) := (others => '0');
    variable b395 : boolean := false;
    variable r394 : std_logic_vector(0 to 17) := (others => '0');
    variable r393 : std_logic_vector(0 to 18) := (others => '0');
    variable b392 : boolean := false;
    variable b391 : boolean := false;
    variable b390 : boolean := false;
    variable r389 : std_logic_vector(0 to 8) := (others => '0');
    variable r388 : std_logic_vector(0 to 8) := (others => '0');
    variable b387 : boolean := false;
    variable r386 : std_logic_vector(0 to 35) := (others => '0');
    variable r385 : std_logic_vector(0 to 17) := (others => '0');
    variable b384 : boolean := false;
    variable b383 : boolean := false;
    variable b382 : boolean := false;
    variable b381 : boolean := false;
    variable r380 : std_logic_vector(0 to 0) := (others => '0');
    variable r379 : std_logic_vector(0 to 8) := (others => '0');
    variable r378 : std_logic_vector(0 to 8) := (others => '0');
    variable b377 : boolean := false;
    variable r376 : std_logic_vector(0 to 17) := (others => '0');
    variable r375 : std_logic_vector(0 to 18) := (others => '0');
    variable r374 : std_logic_vector(0 to 17) := (others => '0');
    variable b373 : boolean := false;
    variable b372 : boolean := false;
    variable b371 : boolean := false;
    variable b370 : boolean := false;
    variable r369 : std_logic_vector(0 to 0) := (others => '0');
    variable r368 : std_logic_vector(0 to 8) := (others => '0');
    variable r367 : std_logic_vector(0 to 8) := (others => '0');
    variable b366 : boolean := false;
    variable r365 : std_logic_vector(0 to 17) := (others => '0');
    variable r364 : std_logic_vector(0 to 18) := (others => '0');
    variable b363 : boolean := false;
    variable b362 : boolean := false;
    variable b361 : boolean := false;
    variable r360 : std_logic_vector(0 to 8) := (others => '0');
    variable r359 : std_logic_vector(0 to 8) := (others => '0');
    variable b358 : boolean := false;
    variable r357 : std_logic_vector(0 to 35) := (others => '0');
    variable r356 : std_logic_vector(0 to 17) := (others => '0');
    variable b355 : boolean := false;
    variable b354 : boolean := false;
    variable b353 : boolean := false;
    variable b352 : boolean := false;
    variable r351 : std_logic_vector(0 to 0) := (others => '0');
    variable r350 : std_logic_vector(0 to 8) := (others => '0');
    variable r349 : std_logic_vector(0 to 8) := (others => '0');
    variable b348 : boolean := false;
    variable r347 : std_logic_vector(0 to 17) := (others => '0');
    variable r346 : std_logic_vector(0 to 7) := (others => '0');
    variable r345 : std_logic_vector(0 to 8) := (others => '0');
    variable r344 : std_logic_vector(0 to 0) := (others => '0');
    variable r343 : std_logic_vector(0 to 18) := (others => '0');
    variable r342 : std_logic_vector(0 to 17) := (others => '0');
    variable b341 : boolean := false;
    variable b340 : boolean := false;
    variable b339 : boolean := false;
    variable b338 : boolean := false;
    variable r337 : std_logic_vector(0 to 0) := (others => '0');
    variable r336 : std_logic_vector(0 to 8) := (others => '0');
    variable r335 : std_logic_vector(0 to 8) := (others => '0');
    variable b334 : boolean := false;
    variable r333 : std_logic_vector(0 to 17) := (others => '0');
    variable r332 : std_logic_vector(0 to 7) := (others => '0');
    variable r331 : std_logic_vector(0 to 8) := (others => '0');
    variable r330 : std_logic_vector(0 to 0) := (others => '0');
    variable r329 : std_logic_vector(0 to 18) := (others => '0');
    variable b328 : boolean := false;
    variable b327 : boolean := false;
    variable b326 : boolean := false;
    variable r325 : std_logic_vector(0 to 8) := (others => '0');
    variable r324 : std_logic_vector(0 to 8) := (others => '0');
    variable b323 : boolean := false;
    variable r322 : std_logic_vector(0 to 35) := (others => '0');
    variable r321 : std_logic_vector(0 to 17) := (others => '0');
    variable b320 : boolean := false;
    variable b319 : boolean := false;
    variable b318 : boolean := false;
    variable b317 : boolean := false;
    variable r316 : std_logic_vector(0 to 0) := (others => '0');
    variable r315 : std_logic_vector(0 to 8) := (others => '0');
    variable r314 : std_logic_vector(0 to 8) := (others => '0');
    variable b313 : boolean := false;
    variable r312 : std_logic_vector(0 to 17) := (others => '0');
    variable r311 : std_logic_vector(0 to 18) := (others => '0');
    variable r310 : std_logic_vector(0 to 17) := (others => '0');
    variable b309 : boolean := false;
    variable b308 : boolean := false;
    variable b307 : boolean := false;
    variable b306 : boolean := false;
    variable r305 : std_logic_vector(0 to 0) := (others => '0');
    variable r304 : std_logic_vector(0 to 8) := (others => '0');
    variable r303 : std_logic_vector(0 to 8) := (others => '0');
    variable b302 : boolean := false;
    variable r301 : std_logic_vector(0 to 17) := (others => '0');
    variable r300 : std_logic_vector(0 to 18) := (others => '0');
    variable b299 : boolean := false;
    variable b298 : boolean := false;
    variable b297 : boolean := false;
    variable r296 : std_logic_vector(0 to 8) := (others => '0');
    variable r295 : std_logic_vector(0 to 8) := (others => '0');
    variable b294 : boolean := false;
    variable r293 : std_logic_vector(0 to 35) := (others => '0');
    variable r292 : std_logic_vector(0 to 17) := (others => '0');
    variable b291 : boolean := false;
    variable b290 : boolean := false;
    variable b289 : boolean := false;
    variable b288 : boolean := false;
    variable r287 : std_logic_vector(0 to 0) := (others => '0');
    variable r286 : std_logic_vector(0 to 8) := (others => '0');
    variable r285 : std_logic_vector(0 to 8) := (others => '0');
    variable b284 : boolean := false;
    variable r283 : std_logic_vector(0 to 17) := (others => '0');
    variable r282 : std_logic_vector(0 to 18) := (others => '0');
    variable r281 : std_logic_vector(0 to 17) := (others => '0');
    variable b280 : boolean := false;
    variable b279 : boolean := false;
    variable b278 : boolean := false;
    variable b277 : boolean := false;
    variable r276 : std_logic_vector(0 to 0) := (others => '0');
    variable r275 : std_logic_vector(0 to 8) := (others => '0');
    variable r274 : std_logic_vector(0 to 8) := (others => '0');
    variable b273 : boolean := false;
    variable r272 : std_logic_vector(0 to 17) := (others => '0');
    variable r271 : std_logic_vector(0 to 18) := (others => '0');
    variable b270 : boolean := false;
    variable b269 : boolean := false;
    variable b268 : boolean := false;
    variable r267 : std_logic_vector(0 to 8) := (others => '0');
    variable r266 : std_logic_vector(0 to 8) := (others => '0');
    variable b265 : boolean := false;
    variable r264 : std_logic_vector(0 to 35) := (others => '0');
    variable r263 : std_logic_vector(0 to 17) := (others => '0');
    variable b262 : boolean := false;
    variable b261 : boolean := false;
    variable b260 : boolean := false;
    variable b259 : boolean := false;
    variable r258 : std_logic_vector(0 to 0) := (others => '0');
    variable r257 : std_logic_vector(0 to 8) := (others => '0');
    variable r256 : std_logic_vector(0 to 8) := (others => '0');
    variable b255 : boolean := false;
    variable r254 : std_logic_vector(0 to 17) := (others => '0');
    variable r253 : std_logic_vector(0 to 18) := (others => '0');
    variable r252 : std_logic_vector(0 to 17) := (others => '0');
    variable b251 : boolean := false;
    variable b250 : boolean := false;
    variable b249 : boolean := false;
    variable b248 : boolean := false;
    variable r247 : std_logic_vector(0 to 0) := (others => '0');
    variable r246 : std_logic_vector(0 to 8) := (others => '0');
    variable r245 : std_logic_vector(0 to 8) := (others => '0');
    variable b244 : boolean := false;
    variable r243 : std_logic_vector(0 to 17) := (others => '0');
    variable r242 : std_logic_vector(0 to 18) := (others => '0');
    variable b241 : boolean := false;
    variable b240 : boolean := false;
    variable b239 : boolean := false;
    variable r238 : std_logic_vector(0 to 8) := (others => '0');
    variable r237 : std_logic_vector(0 to 8) := (others => '0');
    variable b236 : boolean := false;
    variable r235 : std_logic_vector(0 to 35) := (others => '0');
    variable r234 : std_logic_vector(0 to 17) := (others => '0');
    variable b233 : boolean := false;
    variable b232 : boolean := false;
    variable b231 : boolean := false;
    variable b230 : boolean := false;
    variable r229 : std_logic_vector(0 to 0) := (others => '0');
    variable r228 : std_logic_vector(0 to 8) := (others => '0');
    variable r227 : std_logic_vector(0 to 8) := (others => '0');
    variable b226 : boolean := false;
    variable r225 : std_logic_vector(0 to 17) := (others => '0');
    variable r224 : std_logic_vector(0 to 18) := (others => '0');
    variable r223 : std_logic_vector(0 to 17) := (others => '0');
    variable b222 : boolean := false;
    variable b221 : boolean := false;
    variable b220 : boolean := false;
    variable b219 : boolean := false;
    variable r218 : std_logic_vector(0 to 0) := (others => '0');
    variable r217 : std_logic_vector(0 to 8) := (others => '0');
    variable r216 : std_logic_vector(0 to 8) := (others => '0');
    variable b215 : boolean := false;
    variable r214 : std_logic_vector(0 to 17) := (others => '0');
    variable r213 : std_logic_vector(0 to 18) := (others => '0');
    variable b212 : boolean := false;
    variable b211 : boolean := false;
    variable b210 : boolean := false;
    variable r209 : std_logic_vector(0 to 8) := (others => '0');
    variable r208 : std_logic_vector(0 to 8) := (others => '0');
    variable b207 : boolean := false;
    variable r206 : std_logic_vector(0 to 35) := (others => '0');
    variable r205 : std_logic_vector(0 to 17) := (others => '0');
    variable b204 : boolean := false;
    variable b203 : boolean := false;
    variable b202 : boolean := false;
    variable b201 : boolean := false;
    variable r200 : std_logic_vector(0 to 0) := (others => '0');
    variable r199 : std_logic_vector(0 to 8) := (others => '0');
    variable r198 : std_logic_vector(0 to 8) := (others => '0');
    variable b197 : boolean := false;
    variable r196 : std_logic_vector(0 to 17) := (others => '0');
    variable r195 : std_logic_vector(0 to 7) := (others => '0');
    variable r194 : std_logic_vector(0 to 8) := (others => '0');
    variable r193 : std_logic_vector(0 to 0) := (others => '0');
    variable r192 : std_logic_vector(0 to 18) := (others => '0');
    variable r191 : std_logic_vector(0 to 17) := (others => '0');
    variable b190 : boolean := false;
    variable b189 : boolean := false;
    variable b188 : boolean := false;
    variable b187 : boolean := false;
    variable r186 : std_logic_vector(0 to 0) := (others => '0');
    variable r185 : std_logic_vector(0 to 8) := (others => '0');
    variable r184 : std_logic_vector(0 to 8) := (others => '0');
    variable b183 : boolean := false;
    variable r182 : std_logic_vector(0 to 17) := (others => '0');
    variable r181 : std_logic_vector(0 to 7) := (others => '0');
    variable r180 : std_logic_vector(0 to 8) := (others => '0');
    variable r179 : std_logic_vector(0 to 0) := (others => '0');
    variable r178 : std_logic_vector(0 to 18) := (others => '0');
    variable b177 : boolean := false;
    variable b176 : boolean := false;
    variable b175 : boolean := false;
    variable r174 : std_logic_vector(0 to 8) := (others => '0');
    variable r173 : std_logic_vector(0 to 8) := (others => '0');
    variable b172 : boolean := false;
    variable r171 : std_logic_vector(0 to 35) := (others => '0');
    variable r170 : std_logic_vector(0 to 17) := (others => '0');
    variable b169 : boolean := false;
    variable b168 : boolean := false;
    variable b167 : boolean := false;
    variable b166 : boolean := false;
    variable r165 : std_logic_vector(0 to 0) := (others => '0');
    variable r164 : std_logic_vector(0 to 8) := (others => '0');
    variable r163 : std_logic_vector(0 to 8) := (others => '0');
    variable b162 : boolean := false;
    variable r161 : std_logic_vector(0 to 17) := (others => '0');
    variable r160 : std_logic_vector(0 to 18) := (others => '0');
    variable r159 : std_logic_vector(0 to 17) := (others => '0');
    variable b158 : boolean := false;
    variable b157 : boolean := false;
    variable b156 : boolean := false;
    variable b155 : boolean := false;
    variable r154 : std_logic_vector(0 to 0) := (others => '0');
    variable r153 : std_logic_vector(0 to 8) := (others => '0');
    variable r152 : std_logic_vector(0 to 8) := (others => '0');
    variable b151 : boolean := false;
    variable r150 : std_logic_vector(0 to 17) := (others => '0');
    variable r149 : std_logic_vector(0 to 18) := (others => '0');
    variable b148 : boolean := false;
    variable b147 : boolean := false;
    variable b146 : boolean := false;
    variable r145 : std_logic_vector(0 to 8) := (others => '0');
    variable r144 : std_logic_vector(0 to 8) := (others => '0');
    variable b143 : boolean := false;
    variable r142 : std_logic_vector(0 to 35) := (others => '0');
    variable r141 : std_logic_vector(0 to 17) := (others => '0');
    variable b140 : boolean := false;
    variable b139 : boolean := false;
    variable b138 : boolean := false;
    variable b137 : boolean := false;
    variable r136 : std_logic_vector(0 to 0) := (others => '0');
    variable r135 : std_logic_vector(0 to 8) := (others => '0');
    variable r134 : std_logic_vector(0 to 8) := (others => '0');
    variable b133 : boolean := false;
    variable r132 : std_logic_vector(0 to 17) := (others => '0');
    variable r131 : std_logic_vector(0 to 18) := (others => '0');
    variable r130 : std_logic_vector(0 to 17) := (others => '0');
    variable b129 : boolean := false;
    variable b128 : boolean := false;
    variable b127 : boolean := false;
    variable b126 : boolean := false;
    variable r125 : std_logic_vector(0 to 0) := (others => '0');
    variable r124 : std_logic_vector(0 to 8) := (others => '0');
    variable r123 : std_logic_vector(0 to 8) := (others => '0');
    variable b122 : boolean := false;
    variable r121 : std_logic_vector(0 to 17) := (others => '0');
    variable r120 : std_logic_vector(0 to 18) := (others => '0');
    variable b119 : boolean := false;
    variable b118 : boolean := false;
    variable b117 : boolean := false;
    variable r116 : std_logic_vector(0 to 8) := (others => '0');
    variable r115 : std_logic_vector(0 to 8) := (others => '0');
    variable b114 : boolean := false;
    variable r113 : std_logic_vector(0 to 35) := (others => '0');
    variable r112 : std_logic_vector(0 to 17) := (others => '0');
    variable b111 : boolean := false;
    variable b110 : boolean := false;
    variable b109 : boolean := false;
    variable b108 : boolean := false;
    variable r107 : std_logic_vector(0 to 0) := (others => '0');
    variable r106 : std_logic_vector(0 to 8) := (others => '0');
    variable r105 : std_logic_vector(0 to 8) := (others => '0');
    variable b104 : boolean := false;
    variable r103 : std_logic_vector(0 to 17) := (others => '0');
    variable r102 : std_logic_vector(0 to 7) := (others => '0');
    variable r101 : std_logic_vector(0 to 8) := (others => '0');
    variable r100 : std_logic_vector(0 to 0) := (others => '0');
    variable r99 : std_logic_vector(0 to 18) := (others => '0');
    variable r98 : std_logic_vector(0 to 17) := (others => '0');
    variable b97 : boolean := false;
    variable b96 : boolean := false;
    variable b95 : boolean := false;
    variable b94 : boolean := false;
    variable r93 : std_logic_vector(0 to 0) := (others => '0');
    variable r92 : std_logic_vector(0 to 8) := (others => '0');
    variable r91 : std_logic_vector(0 to 8) := (others => '0');
    variable b90 : boolean := false;
    variable r89 : std_logic_vector(0 to 17) := (others => '0');
    variable r88 : std_logic_vector(0 to 7) := (others => '0');
    variable r87 : std_logic_vector(0 to 8) := (others => '0');
    variable r86 : std_logic_vector(0 to 0) := (others => '0');
    variable r85 : std_logic_vector(0 to 18) := (others => '0');
    variable b84 : boolean := false;
    variable b83 : boolean := false;
    variable b82 : boolean := false;
    variable b81 : boolean := false;
    variable b80 : boolean := false;
    variable b79 : boolean := false;
    variable b78 : boolean := false;
    variable b77 : boolean := false;
    variable b76 : boolean := false;
    variable b75 : boolean := false;
    variable b74 : boolean := false;
    variable b73 : boolean := false;
    variable b72 : boolean := false;
    variable b71 : boolean := false;
    variable b70 : boolean := false;
    variable b69 : boolean := false;
    variable b68 : boolean := false;
    variable b67 : boolean := false;
    variable r66 : std_logic_vector(0 to 0) := (others => '0');
    variable r65 : std_logic_vector(0 to 0) := (others => '0');
    variable r64 : std_logic_vector(0 to 0) := (others => '0');
    variable r63 : std_logic_vector(0 to 0) := (others => '0');
    variable r62 : std_logic_vector(0 to 0) := (others => '0');
    variable r61 : std_logic_vector(0 to 0) := (others => '0');
    variable r60 : std_logic_vector(0 to 0) := (others => '0');
    variable r59 : std_logic_vector(0 to 0) := (others => '0');
    variable r58 : std_logic_vector(0 to 0) := (others => '0');
    variable r57 : std_logic_vector(0 to 0) := (others => '0');
    variable r56 : std_logic_vector(0 to 0) := (others => '0');
    variable r55 : std_logic_vector(0 to 0) := (others => '0');
    variable r54 : std_logic_vector(0 to 0) := (others => '0');
    variable r53 : std_logic_vector(0 to 0) := (others => '0');
    variable r52 : std_logic_vector(0 to 0) := (others => '0');
    variable r51 : std_logic_vector(0 to 0) := (others => '0');
    variable b50 : boolean := false;
    variable b49 : boolean := false;
    variable b48 : boolean := false;
    variable b47 : boolean := false;
    variable b46 : boolean := false;
    variable b45 : boolean := false;
    variable r44 : std_logic_vector(0 to 8) := (others => '0');
    variable r43 : std_logic_vector(0 to 8) := (others => '0');
    variable r42 : std_logic_vector(0 to 8) := (others => '0');
    variable r41 : std_logic_vector(0 to 8) := (others => '0');
    variable b40 : boolean := false;
    variable r39 : std_logic_vector(0 to 15) := (others => '0');
    variable r38 : std_logic_vector(0 to 35) := (others => '0');
    variable b37 : boolean := false;
    variable r36 : std_logic_vector(0 to 35) := (others => '0');
    variable r35 : std_logic_vector(0 to 51) := (others => '0');
  begin
    null;
    null;
    null;
    null;
    r35 := (r33 & r34);
    b37 := true;
    r38 := r35(0 to 35);
    r39 := r35(36 to 51);
    b40 := true;
    r41 := r38(0 to 8);
    r42 := r38(9 to 17);
    r43 := r38(18 to 26);
    r44 := r38(27 to 35);
    b45 := true;
    b46 := true;
    b47 := true;
    b48 := true;
    b49 := (b40 AND (b45 AND (b46 AND (b47 AND b48))));
    b50 := true;
    r51 := r39(0 to 0);
    r52 := r39(1 to 1);
    r53 := r39(2 to 2);
    r54 := r39(3 to 3);
    r55 := r39(4 to 4);
    r56 := r39(5 to 5);
    r57 := r39(6 to 6);
    r58 := r39(7 to 7);
    r59 := r39(8 to 8);
    r60 := r39(9 to 9);
    r61 := r39(10 to 10);
    r62 := r39(11 to 11);
    r63 := r39(12 to 12);
    r64 := r39(13 to 13);
    r65 := r39(14 to 14);
    r66 := r39(15 to 15);
    b67 := true;
    b68 := true;
    b69 := true;
    b70 := true;
    b71 := true;
    b72 := true;
    b73 := true;
    b74 := true;
    b75 := true;
    b76 := true;
    b77 := true;
    b78 := true;
    b79 := true;
    b80 := true;
    b81 := true;
    b82 := true;
    b83 := (b50 AND (b67 AND (b68 AND (b69 AND (b70 AND (b71 AND (b72 AND (b73 AND (b74 AND (b75 AND (b76 AND (b77 AND (b78 AND (b79 AND (b80 AND (b81 AND b82))))))))))))))));
    b84 := (b37 AND (b49 AND b83));
    null;
    null;
    null;
    r86 := "0";
    r88 := "00000000";
    r87 := (r86 & r88);
    null;
    r85 := (r44 & r87 & r63);
    b90 := true;
    r91 := r85(0 to 8);
    r92 := r85(9 to 17);
    r93 := r85(18 to 18);
    b94 := true;
    b95 := true;
    b96 := ("1" = r93(0 to 0));
    b97 := (b90 AND (b94 AND (b95 AND b96)));
    if b97 then
      null;
      null;
      null;
      null;
      r98 := (r91 & r91);
      r89 := r98;
     else 
      null;
      null;
      null;
      r100 := "0";
      r102 := "00000000";
      r101 := (r100 & r102);
      null;
      r99 := (r44 & r101 & r63);
      b104 := true;
      r105 := r99(0 to 8);
      r106 := r99(9 to 17);
      r107 := r99(18 to 18);
      b108 := true;
      b109 := true;
      b110 := ("0" = r107(0 to 0));
      b111 := (b104 AND (b108 AND (b109 AND b110)));
      null;
      null;
      null;
      null;
      r112 := (r105 & r106);
      r103 := r112;end if;
    b114 := true;
    r115 := r89(0 to 8);
    r116 := r89(9 to 17);
    b117 := true;
    b118 := true;
    b119 := (b114 AND (b117 AND b118));
    null;
    null;
    null;
    null;
    null;
    r120 := (r43 & r116 & r59);
    b122 := true;
    r123 := r120(0 to 8);
    r124 := r120(9 to 17);
    r125 := r120(18 to 18);
    b126 := true;
    b127 := true;
    b128 := ("1" = r125(0 to 0));
    b129 := (b122 AND (b126 AND (b127 AND b128)));
    if b129 then
      null;
      null;
      null;
      null;
      r130 := (r123 & r123);
      r121 := r130;
     else 
      null;
      null;
      null;
      null;
      null;
      r131 := (r43 & r116 & r59);
      b133 := true;
      r134 := r131(0 to 8);
      r135 := r131(9 to 17);
      r136 := r131(18 to 18);
      b137 := true;
      b138 := true;
      b139 := ("0" = r136(0 to 0));
      b140 := (b133 AND (b137 AND (b138 AND b139)));
      null;
      null;
      null;
      null;
      r141 := (r134 & r135);
      r132 := r141;end if;
    b143 := true;
    r144 := r121(0 to 8);
    r145 := r121(9 to 17);
    b146 := true;
    b147 := true;
    b148 := (b143 AND (b146 AND b147));
    null;
    null;
    null;
    null;
    null;
    r149 := (r42 & r145 & r55);
    b151 := true;
    r152 := r149(0 to 8);
    r153 := r149(9 to 17);
    r154 := r149(18 to 18);
    b155 := true;
    b156 := true;
    b157 := ("1" = r154(0 to 0));
    b158 := (b151 AND (b155 AND (b156 AND b157)));
    if b158 then
      null;
      null;
      null;
      null;
      r159 := (r152 & r152);
      r150 := r159;
     else 
      null;
      null;
      null;
      null;
      null;
      r160 := (r42 & r145 & r55);
      b162 := true;
      r163 := r160(0 to 8);
      r164 := r160(9 to 17);
      r165 := r160(18 to 18);
      b166 := true;
      b167 := true;
      b168 := ("0" = r165(0 to 0));
      b169 := (b162 AND (b166 AND (b167 AND b168)));
      null;
      null;
      null;
      null;
      r170 := (r163 & r164);
      r161 := r170;end if;
    b172 := true;
    r173 := r150(0 to 8);
    r174 := r150(9 to 17);
    b175 := true;
    b176 := true;
    b177 := (b172 AND (b175 AND b176));
    null;
    null;
    null;
    r179 := "0";
    r181 := "00000000";
    r180 := (r179 & r181);
    null;
    r178 := (r115 & r180 & r64);
    b183 := true;
    r184 := r178(0 to 8);
    r185 := r178(9 to 17);
    r186 := r178(18 to 18);
    b187 := true;
    b188 := true;
    b189 := ("1" = r186(0 to 0));
    b190 := (b183 AND (b187 AND (b188 AND b189)));
    if b190 then
      null;
      null;
      null;
      null;
      r191 := (r184 & r184);
      r182 := r191;
     else 
      null;
      null;
      null;
      r193 := "0";
      r195 := "00000000";
      r194 := (r193 & r195);
      null;
      r192 := (r115 & r194 & r64);
      b197 := true;
      r198 := r192(0 to 8);
      r199 := r192(9 to 17);
      r200 := r192(18 to 18);
      b201 := true;
      b202 := true;
      b203 := ("0" = r200(0 to 0));
      b204 := (b197 AND (b201 AND (b202 AND b203)));
      null;
      null;
      null;
      null;
      r205 := (r198 & r199);
      r196 := r205;end if;
    b207 := true;
    r208 := r182(0 to 8);
    r209 := r182(9 to 17);
    b210 := true;
    b211 := true;
    b212 := (b207 AND (b210 AND b211));
    null;
    null;
    null;
    null;
    null;
    r213 := (r144 & r209 & r60);
    b215 := true;
    r216 := r213(0 to 8);
    r217 := r213(9 to 17);
    r218 := r213(18 to 18);
    b219 := true;
    b220 := true;
    b221 := ("1" = r218(0 to 0));
    b222 := (b215 AND (b219 AND (b220 AND b221)));
    if b222 then
      null;
      null;
      null;
      null;
      r223 := (r216 & r216);
      r214 := r223;
     else 
      null;
      null;
      null;
      null;
      null;
      r224 := (r144 & r209 & r60);
      b226 := true;
      r227 := r224(0 to 8);
      r228 := r224(9 to 17);
      r229 := r224(18 to 18);
      b230 := true;
      b231 := true;
      b232 := ("0" = r229(0 to 0));
      b233 := (b226 AND (b230 AND (b231 AND b232)));
      null;
      null;
      null;
      null;
      r234 := (r227 & r228);
      r225 := r234;end if;
    b236 := true;
    r237 := r214(0 to 8);
    r238 := r214(9 to 17);
    b239 := true;
    b240 := true;
    b241 := (b236 AND (b239 AND b240));
    null;
    null;
    null;
    null;
    null;
    r242 := (r173 & r238 & r56);
    b244 := true;
    r245 := r242(0 to 8);
    r246 := r242(9 to 17);
    r247 := r242(18 to 18);
    b248 := true;
    b249 := true;
    b250 := ("1" = r247(0 to 0));
    b251 := (b244 AND (b248 AND (b249 AND b250)));
    if b251 then
      null;
      null;
      null;
      null;
      r252 := (r245 & r245);
      r243 := r252;
     else 
      null;
      null;
      null;
      null;
      null;
      r253 := (r173 & r238 & r56);
      b255 := true;
      r256 := r253(0 to 8);
      r257 := r253(9 to 17);
      r258 := r253(18 to 18);
      b259 := true;
      b260 := true;
      b261 := ("0" = r258(0 to 0));
      b262 := (b255 AND (b259 AND (b260 AND b261)));
      null;
      null;
      null;
      null;
      r263 := (r256 & r257);
      r254 := r263;end if;
    b265 := true;
    r266 := r243(0 to 8);
    r267 := r243(9 to 17);
    b268 := true;
    b269 := true;
    b270 := (b265 AND (b268 AND b269));
    null;
    null;
    null;
    null;
    null;
    r271 := (r41 & r174 & r51);
    b273 := true;
    r274 := r271(0 to 8);
    r275 := r271(9 to 17);
    r276 := r271(18 to 18);
    b277 := true;
    b278 := true;
    b279 := ("1" = r276(0 to 0));
    b280 := (b273 AND (b277 AND (b278 AND b279)));
    if b280 then
      null;
      null;
      null;
      null;
      r281 := (r274 & r274);
      r272 := r281;
     else 
      null;
      null;
      null;
      null;
      null;
      r282 := (r41 & r174 & r51);
      b284 := true;
      r285 := r282(0 to 8);
      r286 := r282(9 to 17);
      r287 := r282(18 to 18);
      b288 := true;
      b289 := true;
      b290 := ("0" = r287(0 to 0));
      b291 := (b284 AND (b288 AND (b289 AND b290)));
      null;
      null;
      null;
      null;
      r292 := (r285 & r286);
      r283 := r292;end if;
    b294 := true;
    r295 := r272(0 to 8);
    r296 := r272(9 to 17);
    b297 := true;
    b298 := true;
    b299 := (b294 AND (b297 AND b298));
    null;
    null;
    null;
    null;
    null;
    r300 := (r295 & r267 & r52);
    b302 := true;
    r303 := r300(0 to 8);
    r304 := r300(9 to 17);
    r305 := r300(18 to 18);
    b306 := true;
    b307 := true;
    b308 := ("1" = r305(0 to 0));
    b309 := (b302 AND (b306 AND (b307 AND b308)));
    if b309 then
      null;
      null;
      null;
      null;
      r310 := (r303 & r303);
      r301 := r310;
     else 
      null;
      null;
      null;
      null;
      null;
      r311 := (r295 & r267 & r52);
      b313 := true;
      r314 := r311(0 to 8);
      r315 := r311(9 to 17);
      r316 := r311(18 to 18);
      b317 := true;
      b318 := true;
      b319 := ("0" = r316(0 to 0));
      b320 := (b313 AND (b317 AND (b318 AND b319)));
      null;
      null;
      null;
      null;
      r321 := (r314 & r315);
      r312 := r321;end if;
    b323 := true;
    r324 := r301(0 to 8);
    r325 := r301(9 to 17);
    b326 := true;
    b327 := true;
    b328 := (b323 AND (b326 AND b327));
    null;
    null;
    null;
    r330 := "0";
    r332 := "00000000";
    r331 := (r330 & r332);
    null;
    r329 := (r208 & r331 & r65);
    b334 := true;
    r335 := r329(0 to 8);
    r336 := r329(9 to 17);
    r337 := r329(18 to 18);
    b338 := true;
    b339 := true;
    b340 := ("1" = r337(0 to 0));
    b341 := (b334 AND (b338 AND (b339 AND b340)));
    if b341 then
      null;
      null;
      null;
      null;
      r342 := (r335 & r335);
      r333 := r342;
     else 
      null;
      null;
      null;
      r344 := "0";
      r346 := "00000000";
      r345 := (r344 & r346);
      null;
      r343 := (r208 & r345 & r65);
      b348 := true;
      r349 := r343(0 to 8);
      r350 := r343(9 to 17);
      r351 := r343(18 to 18);
      b352 := true;
      b353 := true;
      b354 := ("0" = r351(0 to 0));
      b355 := (b348 AND (b352 AND (b353 AND b354)));
      null;
      null;
      null;
      null;
      r356 := (r349 & r350);
      r347 := r356;end if;
    b358 := true;
    r359 := r333(0 to 8);
    r360 := r333(9 to 17);
    b361 := true;
    b362 := true;
    b363 := (b358 AND (b361 AND b362));
    null;
    null;
    null;
    null;
    null;
    r364 := (r237 & r360 & r61);
    b366 := true;
    r367 := r364(0 to 8);
    r368 := r364(9 to 17);
    r369 := r364(18 to 18);
    b370 := true;
    b371 := true;
    b372 := ("1" = r369(0 to 0));
    b373 := (b366 AND (b370 AND (b371 AND b372)));
    if b373 then
      null;
      null;
      null;
      null;
      r374 := (r367 & r367);
      r365 := r374;
     else 
      null;
      null;
      null;
      null;
      null;
      r375 := (r237 & r360 & r61);
      b377 := true;
      r378 := r375(0 to 8);
      r379 := r375(9 to 17);
      r380 := r375(18 to 18);
      b381 := true;
      b382 := true;
      b383 := ("0" = r380(0 to 0));
      b384 := (b377 AND (b381 AND (b382 AND b383)));
      null;
      null;
      null;
      null;
      r385 := (r378 & r379);
      r376 := r385;end if;
    b387 := true;
    r388 := r365(0 to 8);
    r389 := r365(9 to 17);
    b390 := true;
    b391 := true;
    b392 := (b387 AND (b390 AND b391));
    null;
    null;
    null;
    null;
    null;
    r393 := (r266 & r389 & r57);
    b395 := true;
    r396 := r393(0 to 8);
    r397 := r393(9 to 17);
    r398 := r393(18 to 18);
    b399 := true;
    b400 := true;
    b401 := ("1" = r398(0 to 0));
    b402 := (b395 AND (b399 AND (b400 AND b401)));
    if b402 then
      null;
      null;
      null;
      null;
      r403 := (r396 & r396);
      r394 := r403;
     else 
      null;
      null;
      null;
      null;
      null;
      r404 := (r266 & r389 & r57);
      b406 := true;
      r407 := r404(0 to 8);
      r408 := r404(9 to 17);
      r409 := r404(18 to 18);
      b410 := true;
      b411 := true;
      b412 := ("0" = r409(0 to 0));
      b413 := (b406 AND (b410 AND (b411 AND b412)));
      null;
      null;
      null;
      null;
      r414 := (r407 & r408);
      r405 := r414;end if;
    b416 := true;
    r417 := r394(0 to 8);
    r418 := r394(9 to 17);
    b419 := true;
    b420 := true;
    b421 := (b416 AND (b419 AND b420));
    null;
    null;
    null;
    null;
    null;
    r422 := (r324 & r418 & r53);
    b424 := true;
    r425 := r422(0 to 8);
    r426 := r422(9 to 17);
    r427 := r422(18 to 18);
    b428 := true;
    b429 := true;
    b430 := ("1" = r427(0 to 0));
    b431 := (b424 AND (b428 AND (b429 AND b430)));
    if b431 then
      null;
      null;
      null;
      null;
      r432 := (r425 & r425);
      r423 := r432;
     else 
      null;
      null;
      null;
      null;
      null;
      r433 := (r324 & r418 & r53);
      b435 := true;
      r436 := r433(0 to 8);
      r437 := r433(9 to 17);
      r438 := r433(18 to 18);
      b439 := true;
      b440 := true;
      b441 := ("0" = r438(0 to 0));
      b442 := (b435 AND (b439 AND (b440 AND b441)));
      null;
      null;
      null;
      null;
      r443 := (r436 & r437);
      r434 := r443;end if;
    b445 := true;
    r446 := r423(0 to 8);
    r447 := r423(9 to 17);
    b448 := true;
    b449 := true;
    b450 := (b445 AND (b448 AND b449));
    null;
    null;
    null;
    r452 := "0";
    r454 := "00000000";
    r453 := (r452 & r454);
    null;
    r451 := (r359 & r453 & r66);
    b456 := true;
    r457 := r451(0 to 8);
    r458 := r451(9 to 17);
    r459 := r451(18 to 18);
    b460 := true;
    b461 := true;
    b462 := ("1" = r459(0 to 0));
    b463 := (b456 AND (b460 AND (b461 AND b462)));
    if b463 then
      null;
      null;
      null;
      null;
      r464 := (r457 & r457);
      r455 := r464;
     else 
      null;
      null;
      null;
      r466 := "0";
      r468 := "00000000";
      r467 := (r466 & r468);
      null;
      r465 := (r359 & r467 & r66);
      b470 := true;
      r471 := r465(0 to 8);
      r472 := r465(9 to 17);
      r473 := r465(18 to 18);
      b474 := true;
      b475 := true;
      b476 := ("0" = r473(0 to 0));
      b477 := (b470 AND (b474 AND (b475 AND b476)));
      null;
      null;
      null;
      null;
      r478 := (r471 & r472);
      r469 := r478;end if;
    b480 := true;
    r481 := r455(0 to 8);
    r482 := r455(9 to 17);
    b483 := true;
    b484 := true;
    b485 := (b480 AND (b483 AND b484));
    null;
    null;
    null;
    null;
    null;
    r486 := (r388 & r482 & r62);
    b488 := true;
    r489 := r486(0 to 8);
    r490 := r486(9 to 17);
    r491 := r486(18 to 18);
    b492 := true;
    b493 := true;
    b494 := ("1" = r491(0 to 0));
    b495 := (b488 AND (b492 AND (b493 AND b494)));
    if b495 then
      null;
      null;
      null;
      null;
      r496 := (r489 & r489);
      r487 := r496;
     else 
      null;
      null;
      null;
      null;
      null;
      r497 := (r388 & r482 & r62);
      b499 := true;
      r500 := r497(0 to 8);
      r501 := r497(9 to 17);
      r502 := r497(18 to 18);
      b503 := true;
      b504 := true;
      b505 := ("0" = r502(0 to 0));
      b506 := (b499 AND (b503 AND (b504 AND b505)));
      null;
      null;
      null;
      null;
      r507 := (r500 & r501);
      r498 := r507;end if;
    b509 := true;
    r510 := r487(0 to 8);
    r511 := r487(9 to 17);
    b512 := true;
    b513 := true;
    b514 := (b509 AND (b512 AND b513));
    null;
    null;
    null;
    null;
    null;
    r515 := (r417 & r511 & r58);
    b517 := true;
    r518 := r515(0 to 8);
    r519 := r515(9 to 17);
    r520 := r515(18 to 18);
    b521 := true;
    b522 := true;
    b523 := ("1" = r520(0 to 0));
    b524 := (b517 AND (b521 AND (b522 AND b523)));
    if b524 then
      null;
      null;
      null;
      null;
      r525 := (r518 & r518);
      r516 := r525;
     else 
      null;
      null;
      null;
      null;
      null;
      r526 := (r417 & r511 & r58);
      b528 := true;
      r529 := r526(0 to 8);
      r530 := r526(9 to 17);
      r531 := r526(18 to 18);
      b532 := true;
      b533 := true;
      b534 := ("0" = r531(0 to 0));
      b535 := (b528 AND (b532 AND (b533 AND b534)));
      null;
      null;
      null;
      null;
      r536 := (r529 & r530);
      r527 := r536;end if;
    b538 := true;
    r539 := r516(0 to 8);
    r540 := r516(9 to 17);
    b541 := true;
    b542 := true;
    b543 := (b538 AND (b541 AND b542));
    null;
    null;
    null;
    null;
    null;
    r544 := (r446 & r540 & r54);
    b546 := true;
    r547 := r544(0 to 8);
    r548 := r544(9 to 17);
    r549 := r544(18 to 18);
    b550 := true;
    b551 := true;
    b552 := ("1" = r549(0 to 0));
    b553 := (b546 AND (b550 AND (b551 AND b552)));
    if b553 then
      null;
      null;
      null;
      null;
      r554 := (r547 & r547);
      r545 := r554;
     else 
      null;
      null;
      null;
      null;
      null;
      r555 := (r446 & r540 & r54);
      b557 := true;
      r558 := r555(0 to 8);
      r559 := r555(9 to 17);
      r560 := r555(18 to 18);
      b561 := true;
      b562 := true;
      b563 := ("0" = r560(0 to 0));
      b564 := (b557 AND (b561 AND (b562 AND b563)));
      null;
      null;
      null;
      null;
      r565 := (r558 & r559);
      r556 := r565;end if;
    b567 := true;
    r568 := r545(0 to 8);
    r569 := r545(9 to 17);
    b570 := true;
    b571 := true;
    b572 := (b567 AND (b570 AND b571));
    null;
    null;
    null;
    null;
    null;
    null;
    r573 := (r296 & r325 & r447 & r569);
    r566 := r573;
    r537 := r566;
    r508 := r537;
    r479 := r508;
    r444 := r479;
    r415 := r444;
    r386 := r415;
    r357 := r386;
    r322 := r357;
    r293 := r322;
    r264 := r293;
    r235 := r264;
    r206 := r235;
    r171 := r206;
    r142 := r171;
    r113 := r142;
    r36 := r113;
    return r36;
  end rewire_Maincrossbar_32;
  signal control_flop : control_state := STATE0;
  signal control_flop_next : control_state := STATE0;
  signal input_flop : std_logic_vector(0 to 52) := (others => '0');
  signal goto_L604_flop : boolean := false;
  signal goto_L597_flop : boolean := false;
  signal goto_L581_flop : boolean := false;
  signal goto_L11_flop : boolean := false;
  signal goto_L13_flop : boolean := false;
  signal goto_L585_flop : boolean := false;
  signal goto_L29_flop : boolean := false;
  signal goto_L0_flop : boolean := false;
  signal goto_L605_flop : boolean := false;
  signal r596_flop : std_logic_vector(0 to 52) := (others => '0');
  signal r592_flop : std_logic_vector(0 to 35) := (others => '0');
  signal r591_flop : std_logic_vector(0 to 36) := (others => '0');
  signal r589_flop : std_logic_vector(0 to 0) := (others => '0');
  signal r580_flop : std_logic_vector(0 to 52) := (others => '0');
  signal r576_flop : std_logic_vector(0 to 35) := (others => '0');
  signal r34_flop : std_logic_vector(0 to 15) := (others => '0');
  signal r33_flop : std_logic_vector(0 to 35) := (others => '0');
  signal r30_flop : std_logic_vector(0 to 36) := (others => '0');
  signal r28_flop : std_logic_vector(0 to 0) := (others => '0');
  signal b26_flop : boolean := false;
  signal b24_flop : boolean := false;
  signal b22_flop : boolean := false;
  signal r20_flop : std_logic_vector(0 to 15) := (others => '0');
  signal r18_flop : std_logic_vector(0 to 35) := (others => '0');
  signal b16_flop : boolean := false;
  signal r12_flop : std_logic_vector(0 to 52) := (others => '0');
  signal r10_flop : std_logic_vector(0 to 52) := (others => '0');
  signal r6_flop : std_logic_vector(0 to 35) := (others => '0');
  signal r5_flop : std_logic_vector(0 to 36) := (others => '0');
  signal r3_flop : std_logic_vector(0 to 0) := (others => '0');
  signal goto_L604_flop_next : boolean := false;
  signal goto_L597_flop_next : boolean := false;
  signal goto_L581_flop_next : boolean := false;
  signal goto_L11_flop_next : boolean := false;
  signal goto_L13_flop_next : boolean := false;
  signal goto_L585_flop_next : boolean := false;
  signal goto_L29_flop_next : boolean := false;
  signal goto_L0_flop_next : boolean := false;
  signal goto_L605_flop_next : boolean := false;
  signal r596_flop_next : std_logic_vector(0 to 52) := (others => '0');
  signal r592_flop_next : std_logic_vector(0 to 35) := (others => '0');
  signal r591_flop_next : std_logic_vector(0 to 36) := (others => '0');
  signal r589_flop_next : std_logic_vector(0 to 0) := (others => '0');
  signal r580_flop_next : std_logic_vector(0 to 52) := (others => '0');
  signal r576_flop_next : std_logic_vector(0 to 35) := (others => '0');
  signal r34_flop_next : std_logic_vector(0 to 15) := (others => '0');
  signal r33_flop_next : std_logic_vector(0 to 35) := (others => '0');
  signal r30_flop_next : std_logic_vector(0 to 36) := (others => '0');
  signal r28_flop_next : std_logic_vector(0 to 0) := (others => '0');
  signal b26_flop_next : boolean := false;
  signal b24_flop_next : boolean := false;
  signal b22_flop_next : boolean := false;
  signal r20_flop_next : std_logic_vector(0 to 15) := (others => '0');
  signal r18_flop_next : std_logic_vector(0 to 35) := (others => '0');
  signal b16_flop_next : boolean := false;
  signal r12_flop_next : std_logic_vector(0 to 52) := (others => '0');
  signal r10_flop_next : std_logic_vector(0 to 52) := (others => '0');
  signal r6_flop_next : std_logic_vector(0 to 35) := (others => '0');
  signal r5_flop_next : std_logic_vector(0 to 36) := (others => '0');
  signal r3_flop_next : std_logic_vector(0 to 0) := (others => '0');
begin
  -- Logic loop process.
  process (control_flop,input_flop,goto_L604_flop,goto_L597_flop,goto_L581_flop,goto_L11_flop,goto_L13_flop,goto_L585_flop,goto_L29_flop,goto_L0_flop,goto_L605_flop,r596_flop,r592_flop,r591_flop,r589_flop,r580_flop,r576_flop,r34_flop,r33_flop,r30_flop,r28_flop,b26_flop,b24_flop,b22_flop,r20_flop,r18_flop,b16_flop,r12_flop,r10_flop,r6_flop,r5_flop,r3_flop)
    variable control : control_state;
    variable input_tmp : std_logic_vector(0 to 52);
    variable goto_L604 : boolean := false;
    variable goto_L597 : boolean := false;
    variable goto_L581 : boolean := false;
    variable goto_L11 : boolean := false;
    variable goto_L13 : boolean := false;
    variable goto_L585 : boolean := false;
    variable goto_L29 : boolean := false;
    variable goto_L0 : boolean := false;
    variable goto_L605 : boolean := false;
    variable r596 : std_logic_vector(0 to 52) := (others => '0');
    variable r592 : std_logic_vector(0 to 35) := (others => '0');
    variable r591 : std_logic_vector(0 to 36) := (others => '0');
    variable r589 : std_logic_vector(0 to 0) := (others => '0');
    variable r580 : std_logic_vector(0 to 52) := (others => '0');
    variable r576 : std_logic_vector(0 to 35) := (others => '0');
    variable r34 : std_logic_vector(0 to 15) := (others => '0');
    variable r33 : std_logic_vector(0 to 35) := (others => '0');
    variable r30 : std_logic_vector(0 to 36) := (others => '0');
    variable r28 : std_logic_vector(0 to 0) := (others => '0');
    variable b26 : boolean := false;
    variable b24 : boolean := false;
    variable b22 : boolean := false;
    variable r20 : std_logic_vector(0 to 15) := (others => '0');
    variable r18 : std_logic_vector(0 to 35) := (others => '0');
    variable b16 : boolean := false;
    variable r12 : std_logic_vector(0 to 52) := (others => '0');
    variable r10 : std_logic_vector(0 to 52) := (others => '0');
    variable r6 : std_logic_vector(0 to 35) := (others => '0');
    variable r5 : std_logic_vector(0 to 36) := (others => '0');
    variable r3 : std_logic_vector(0 to 0) := (others => '0');
    variable output_tmp : std_logic_vector(0 to 36);
  begin
    -- Read reg temps.
    control := control_flop;
    input_tmp := input_flop;
    goto_L604 := goto_L604_flop;
    goto_L597 := goto_L597_flop;
    goto_L581 := goto_L581_flop;
    goto_L11 := goto_L11_flop;
    goto_L13 := goto_L13_flop;
    goto_L585 := goto_L585_flop;
    goto_L29 := goto_L29_flop;
    goto_L0 := goto_L0_flop;
    goto_L605 := goto_L605_flop;
    r596 := r596_flop;
    r592 := r592_flop;
    r591 := r591_flop;
    r589 := r589_flop;
    r580 := r580_flop;
    r576 := r576_flop;
    r34 := r34_flop;
    r33 := r33_flop;
    r30 := r30_flop;
    r28 := r28_flop;
    b26 := b26_flop;
    b24 := b24_flop;
    b22 := b22_flop;
    r20 := r20_flop;
    r18 := r18_flop;
    b16 := b16_flop;
    r12 := r12_flop;
    r10 := r10_flop;
    r6 := r6_flop;
    r5 := r5_flop;
    r3 := r3_flop;
    output_tmp := (others => '0');
    -- Loop body.
    goto_L604 := false;
    goto_L597 := false;
    goto_L581 := false;
    goto_L11 := false;
    goto_L13 := false;
    goto_L585 := false;
    goto_L29 := false;
    goto_L0 := false;
    goto_L605 := false;
    null; -- label L604
    -- ENTER
    goto_L0 := (control = STATE0);
    if (NOT goto_L0) then
      goto_L11 := (control = STATE11);
      if (NOT goto_L11) then
        goto_L581 := (control = STATE581);
        if (NOT goto_L581) then
          goto_L597 := (control = STATE597);
          null; -- label L597
          r596 := input_tmp;
          -- got i@215 in r596
          r12 := r596;
          goto_L13 := true;
        end if;
        goto_L13 := goto_L13;
        if (NOT goto_L13) then
          null; -- label L581
          r580 := input_tmp;
          -- got i@214 in r580
          r12 := r580;
          goto_L13 := true;
        end if;
        goto_L13 := goto_L13;
      end if;
      goto_L13 := goto_L13;
      if (NOT goto_L13) then
        null; -- label L11
        r10 := input_tmp;
        -- got i@210 in r10
        r12 := r10;
        goto_L13 := true;
      end if;
      goto_L13 := goto_L13;
      null; -- label L13
      -- Main.dev in
      -- got $5@211 in r12
      b16 := ("0" = r12(0 to 0));
      r18 := r12(1 to 36);
      r20 := r12(37 to 52);
      b22 := true;
      b24 := true;
      b26 := (b16 AND (b22 AND b24));
      goto_L29 := b26;
      if (NOT goto_L29) then
        goto_L585 := (NOT b26);
        null; -- label L585
        -- alt exit (no match)
        -- got $5@211 in r12
        -- final pat
        r589 := "1";
        r592 := "000000000000000000000000000000000000";
        r591 := (r589 & r592);
        output_tmp := r591;
        control := STATE597;
        goto_L605 := true;
      end if;
      goto_L605 := goto_L605;
      if (NOT goto_L605) then
        null; -- label L29
        r28 := "0";
        null;
        -- got m4@212 in r18
        -- got b16@213 in r20
        r576 := rewire_Maincrossbar_32(r18,r20);
        r30 := (r28 & r576);
        output_tmp := r30;
        control := STATE581;
        goto_L605 := true;
      end if;
      goto_L605 := goto_L605;
    end if;
    goto_L605 := goto_L605;
    if (NOT goto_L605) then
      null; -- label L0
      -- START
      -- Main.devcrossbar in
      r3 := "1";
      r6 := "000000000000000000000000000000000000";
      r5 := (r3 & r6);
      output_tmp := r5;
      control := STATE11;
      goto_L605 := true;
    end if;
    goto_L605 := goto_L605;
    null; -- label L605
    -- EXIT
    -- Write back reg temps.
    control_flop_next <= control;
    goto_L604_flop_next <= goto_L604;
    goto_L597_flop_next <= goto_L597;
    goto_L581_flop_next <= goto_L581;
    goto_L11_flop_next <= goto_L11;
    goto_L13_flop_next <= goto_L13;
    goto_L585_flop_next <= goto_L585;
    goto_L29_flop_next <= goto_L29;
    goto_L0_flop_next <= goto_L0;
    goto_L605_flop_next <= goto_L605;
    r596_flop_next <= r596;
    r592_flop_next <= r592;
    r591_flop_next <= r591;
    r589_flop_next <= r589;
    r580_flop_next <= r580;
    r576_flop_next <= r576;
    r34_flop_next <= r34;
    r33_flop_next <= r33;
    r30_flop_next <= r30;
    r28_flop_next <= r28;
    b26_flop_next <= b26;
    b24_flop_next <= b24;
    b22_flop_next <= b22;
    r20_flop_next <= r20;
    r18_flop_next <= r18;
    b16_flop_next <= b16;
    r12_flop_next <= r12;
    r10_flop_next <= r10;
    r6_flop_next <= r6;
    r5_flop_next <= r5;
    r3_flop_next <= r3;
    -- Update output line.
    output <= output_tmp;
  end process;

  -- Flip flop update process.
  process (clk,input,goto_L604_flop_next,goto_L597_flop_next,goto_L581_flop_next,goto_L11_flop_next,goto_L13_flop_next,goto_L585_flop_next,goto_L29_flop_next,goto_L0_flop_next,goto_L605_flop_next,r596_flop_next,r592_flop_next,r591_flop_next,r589_flop_next,r580_flop_next,r576_flop_next,r34_flop_next,r33_flop_next,r30_flop_next,r28_flop_next,b26_flop_next,b24_flop_next,b22_flop_next,r20_flop_next,r18_flop_next,b16_flop_next,r12_flop_next,r10_flop_next,r6_flop_next,r5_flop_next,r3_flop_next)
  begin
    if clk'event and clk='1' then
      input_flop <= input;
      control_flop <= control_flop_next;
      goto_L604_flop <= goto_L604_flop_next;
      goto_L597_flop <= goto_L597_flop_next;
      goto_L581_flop <= goto_L581_flop_next;
      goto_L11_flop <= goto_L11_flop_next;
      goto_L13_flop <= goto_L13_flop_next;
      goto_L585_flop <= goto_L585_flop_next;
      goto_L29_flop <= goto_L29_flop_next;
      goto_L0_flop <= goto_L0_flop_next;
      goto_L605_flop <= goto_L605_flop_next;
      r596_flop <= r596_flop_next;
      r592_flop <= r592_flop_next;
      r591_flop <= r591_flop_next;
      r589_flop <= r589_flop_next;
      r580_flop <= r580_flop_next;
      r576_flop <= r576_flop_next;
      r34_flop <= r34_flop_next;
      r33_flop <= r33_flop_next;
      r30_flop <= r30_flop_next;
      r28_flop <= r28_flop_next;
      b26_flop <= b26_flop_next;
      b24_flop <= b24_flop_next;
      b22_flop <= b22_flop_next;
      r20_flop <= r20_flop_next;
      r18_flop <= r18_flop_next;
      b16_flop <= b16_flop_next;
      r12_flop <= r12_flop_next;
      r10_flop <= r10_flop_next;
      r6_flop <= r6_flop_next;
      r5_flop <= r5_flop_next;
      r3_flop <= r3_flop_next;
    end if;
  end process;

end behavioral;
